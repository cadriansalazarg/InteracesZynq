`timescale 1ns / 1ps

//`define PACKET_SIZE_4096
//`define PACKET_SIZE_2048
`define PACKET_SIZE_1024  //Debe ajustarse al tamaño de paquete que mejor se ajusta, de manera que concuerde con PACKET_SIZE_BITS, o al menos PACKET_SIZE_BITS sea menor o igual que este parámetro
//`define PACKET_SIZE_512
//`define PACKET_SIZE_256

// Descripción de parámetros
// PACKET_SIZE_BITS representa el tamaño del paquete en bits,los valores testeados son 256, 512 y 1024. Sin embargo debería se servir bien hasta 4096
// NUMBER_OF_LANES representa el número de lanes para los que fue configurado el Aurora, solo fue testeado con dos lanes, por lo tanto, solo puede usarse el valor de 1, o el valor de 2
// DATAFILE es un parámetro que permite variar el contenido de la memoria ROM que se encarga de generar el BS_ID en función del valor de RX_UID. Los diferentes archivos de que se deberán de cargar en la ROM deben de llamarse como Memory_Content_X.txt, donde X puede ser 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, de esta manera cambiando este parámetro, se puede usar este bloque en para dferentes FPGAs

module Aurora_to_fifo #(parameter PACKET_SIZE_BITS = 256, parameter NUMBER_OF_LANES = 1, parameter DATAFILE = 1)
(user_clk, reset_TX_RX_Block,  din, wr_en, m_axi_rx_tdata, m_axi_rx_tlast, m_axi_rx_tvalid, full, Error);

    localparam n = 32*NUMBER_OF_LANES; 
    
    localparam S0 = 3'd0, S1 = 3'd1, S2 = 3'd2, S3 = 3'd3, S4 = 3'd4;
	reg [2:0] State, NextState;

    input user_clk, reset_TX_RX_Block;
    input m_axi_rx_tlast, m_axi_rx_tvalid;
    input [(32*NUMBER_OF_LANES)-1:0] m_axi_rx_tdata;
    input full;
    
    output [PACKET_SIZE_BITS-1: 0] din;
    output reg wr_en;
    output reg Error;
    
     
     
    reg full_reg;
    reg [(32*NUMBER_OF_LANES)-1:0] m_axi_rx_tdata_reg;
    reg [(32*NUMBER_OF_LANES)-1:0] m_axi_rx_tdata_reg1;
    wire [7:0] BS_ID;
    
    
    reg m_axi_rx_tvalid_reg, m_axi_rx_tlast_reg;
    wire [PACKET_SIZE_BITS-1: 0] din_reg;
    reg reset_output_register, wr_en_reg, reset_file_register, enable_output_register;
    reg [7:0] Q_seq_counter;
    
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Registro paralelo paralelo
    // Tiene la función de reducir problemas temporales, al evitar rutas combinacionales
    // largas. Por lo tanto, todas las señales de entrada y salida se almacenan
    // en un registro, previo a su salida al exterior
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
    always @(posedge user_clk) begin
        if (reset_TX_RX_Block) begin
            m_axi_rx_tvalid_reg <= 1'b0;
            m_axi_rx_tlast_reg <= 1'b0;
            m_axi_rx_tdata_reg <= 0;
            full_reg <= 0;
            wr_en <= 0;
        end else begin
            m_axi_rx_tvalid_reg <= m_axi_rx_tvalid;
            m_axi_rx_tlast_reg <= m_axi_rx_tlast;
            m_axi_rx_tdata_reg <= m_axi_rx_tdata;
            full_reg <= full;
            wr_en <= wr_en_reg;
        end
    end
    
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Registro paralelo paralelo con enable
    // Es un segundo registro paralelo paralelo que almacena los datos que salen
    // del Aurora por el puesto m_axi_rx_tdata, pero los datos solo se almacenan 
    // si la señal de valid se encuentra en alto.
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
    
    always @(posedge user_clk) begin
		if (reset_TX_RX_Block) begin 
			m_axi_rx_tdata_reg1 <= 0;
		end else if (m_axi_rx_tvalid_reg) begin
			m_axi_rx_tdata_reg1 <= m_axi_rx_tdata_reg;
		end
	end
    
    
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Registro paralelo paralelo
    // Se instancia en un generate un registro paralelo pralelo, que va a almacenar todos
    // los datos que vienen del Aurora, en un paquete. Note que a todos los registros
    // generados por el generate, les ingresa el mismo Data_Input (m_axi_rx_tdata_reg1)
    // pero solo se habilita el enable de uno de ellos por ciclo de reloj, de esta forma
    // se realiza la construcción del paquete.
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
    
    // Declare a temporary loop variable to be used during
    // genaration and won't be available during simulation
    genvar i;
    
    wire [n-1:0] OutputReg [0:((PACKET_SIZE_BITS/n)-1)];
    wire [(PACKET_SIZE_BITS/n)-1: 0] enable;
    
    generate
        for (i = 0; i<(PACKET_SIZE_BITS/n); i = i + 1) begin
            register #(.WIDTH(n) ) u0(
                .clk(user_clk),
                .reset(reset_TX_RX_Block),
                .enable(Enable_Registers[i]),
                .Din(m_axi_rx_tdata_reg1),
                .Dout(din_reg[ (((PACKET_SIZE_BITS)-1)-(i*n)) :  (((PACKET_SIZE_BITS)-n)-(i*n)) ]));
        end
    endgenerate
    
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Contador binario y decodificador para habilitar el enable
    // Se crea un contador binario y un decodificador con registro a la salida para evitar problemas de timing
    // El contador tiene como enable la señal de valid, de esta forma, solo cuando existan datos válidos este podrá contar.
    // La salida del contador se conecta al puerto de entrada del decodificador, de esta forma, con cada flanco de reloj, 
    // se habilitará un registro diferente del banco de registros, almacenando así el dato en diferentes posiciones.
    // Se usa un if_def en función del tamaño del paquete. 
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
    
    
    // *********************************** Counter and decoder in function of packet size ********************************
`ifdef PACKET_SIZE_4096
	reg [6:0] Q_counter;
	reg [127:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				7'd0  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
				7'd1  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
				7'd2  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
				7'd3  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
				7'd4  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
				7'd5  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
				7'd6  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
				7'd7  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
				7'd8  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
				7'd9  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
				7'd10 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
				7'd11 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
				7'd12 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
				7'd13 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
				7'd14 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
				7'd15 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;	
				7'd16 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
				7'd17 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
				7'd18 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
				7'd19 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
				7'd20 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
				7'd21 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
				7'd22 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
				7'd23 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
				7'd24 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
				7'd25 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
				7'd26 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
				7'd27 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
				7'd28 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
				7'd29 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
				7'd30 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
				7'd31 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
				7'd32 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
				7'd33 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
				7'd34 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
				7'd35 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
				7'd36 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
				7'd37 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
				7'd38 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
				7'd39 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
				7'd40 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
				7'd41 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
				7'd42 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
				7'd43 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
				7'd44 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
				7'd45 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
				7'd46 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
				7'd47 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;	
				7'd48 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
				7'd49 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
				7'd50 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
				7'd51 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
				7'd52 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
				7'd53 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
				7'd54 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
				7'd55 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
				7'd56 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
				7'd57 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
				7'd58 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
				7'd59 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
				7'd60 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
				7'd61 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
				7'd62 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
				7'd63 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
				7'd64 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
				7'd65 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
				7'd66 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
				7'd67 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
				7'd68 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
				7'd69 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
				7'd70 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
				7'd71 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
				7'd72 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd73 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd74 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd75 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd76 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd77 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd78 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd79 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;	
				7'd80 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd81 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd82 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd83 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd84 : Enable_Registers <= 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd85 : Enable_Registers <= 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd86 : Enable_Registers <= 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd87 : Enable_Registers <= 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd88 : Enable_Registers <= 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd89 : Enable_Registers <= 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd90 : Enable_Registers <= 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd91 : Enable_Registers <= 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd92 : Enable_Registers <= 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd93 : Enable_Registers <= 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd94 : Enable_Registers <= 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd95 : Enable_Registers <= 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd96 : Enable_Registers <= 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd97 : Enable_Registers <= 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd98 : Enable_Registers <= 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd99 : Enable_Registers <= 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd100: Enable_Registers <= 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd101: Enable_Registers <= 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd102: Enable_Registers <= 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd103: Enable_Registers <= 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd104: Enable_Registers <= 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd105: Enable_Registers <= 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd106: Enable_Registers <= 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd107: Enable_Registers <= 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd108: Enable_Registers <= 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd109: Enable_Registers <= 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd110: Enable_Registers <= 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd111: Enable_Registers <= 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;	
				7'd112: Enable_Registers <= 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd113: Enable_Registers <= 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd114: Enable_Registers <= 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd115: Enable_Registers <= 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd116: Enable_Registers <= 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd117: Enable_Registers <= 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd118: Enable_Registers <= 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd119: Enable_Registers <= 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd120: Enable_Registers <= 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd121: Enable_Registers <= 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd122: Enable_Registers <= 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd123: Enable_Registers <= 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd124: Enable_Registers <= 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd125: Enable_Registers <= 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd126: Enable_Registers <= 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd127: Enable_Registers <= 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_2048
	reg [5:0] Q_counter;
	reg [63:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				6'd0  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
				6'd1  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
				6'd2  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
				6'd3  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
				6'd4  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
				6'd5  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
				6'd6  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
				6'd7  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
				6'd8  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
				6'd9  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000001000000000;
				6'd10 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000010000000000;
				6'd11 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000100000000000;
				6'd12 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000001000000000000;
				6'd13 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000010000000000000;
				6'd14 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000100000000000000;
				6'd15 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000001000000000000000;	
				6'd16 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000010000000000000000;
				6'd17 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000100000000000000000;
				6'd18 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
				6'd19 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000010000000000000000000;
				6'd20 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000100000000000000000000;
				6'd21 : Enable_Registers <= 64'b0000000000000000000000000000000000000000001000000000000000000000;
				6'd22 : Enable_Registers <= 64'b0000000000000000000000000000000000000000010000000000000000000000;
				6'd23 : Enable_Registers <= 64'b0000000000000000000000000000000000000000100000000000000000000000;
				6'd24 : Enable_Registers <= 64'b0000000000000000000000000000000000000001000000000000000000000000;
				6'd25 : Enable_Registers <= 64'b0000000000000000000000000000000000000010000000000000000000000000;
				6'd26 : Enable_Registers <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
				6'd27 : Enable_Registers <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
				6'd28 : Enable_Registers <= 64'b0000000000000000000000000000000000010000000000000000000000000000;
				6'd29 : Enable_Registers <= 64'b0000000000000000000000000000000000100000000000000000000000000000;
				6'd30 : Enable_Registers <= 64'b0000000000000000000000000000000001000000000000000000000000000000;
				6'd31 : Enable_Registers <= 64'b0000000000000000000000000000000010000000000000000000000000000000;
				6'd32 : Enable_Registers <= 64'b0000000000000000000000000000000100000000000000000000000000000000;
				6'd33 : Enable_Registers <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
				6'd34 : Enable_Registers <= 64'b0000000000000000000000000000010000000000000000000000000000000000;
				6'd35 : Enable_Registers <= 64'b0000000000000000000000000000100000000000000000000000000000000000;
				6'd36 : Enable_Registers <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
				6'd37 : Enable_Registers <= 64'b0000000000000000000000000010000000000000000000000000000000000000;
				6'd38 : Enable_Registers <= 64'b0000000000000000000000000100000000000000000000000000000000000000;
				6'd39 : Enable_Registers <= 64'b0000000000000000000000001000000000000000000000000000000000000000;
				6'd40 : Enable_Registers <= 64'b0000000000000000000000010000000000000000000000000000000000000000;
				6'd41 : Enable_Registers <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
				6'd42 : Enable_Registers <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
				6'd43 : Enable_Registers <= 64'b0000000000000000000010000000000000000000000000000000000000000000;
				6'd44 : Enable_Registers <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
				6'd45 : Enable_Registers <= 64'b0000000000000000001000000000000000000000000000000000000000000000;
				6'd46 : Enable_Registers <= 64'b0000000000000000010000000000000000000000000000000000000000000000;
				6'd47 : Enable_Registers <= 64'b0000000000000000100000000000000000000000000000000000000000000000;	
				6'd48 : Enable_Registers <= 64'b0000000000000001000000000000000000000000000000000000000000000000;
				6'd49 : Enable_Registers <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
				6'd50 : Enable_Registers <= 64'b0000000000000100000000000000000000000000000000000000000000000000;
				6'd51 : Enable_Registers <= 64'b0000000000001000000000000000000000000000000000000000000000000000;
				6'd52 : Enable_Registers <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				6'd53 : Enable_Registers <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
				6'd54 : Enable_Registers <= 64'b0000000001000000000000000000000000000000000000000000000000000000;
				6'd55 : Enable_Registers <= 64'b0000000010000000000000000000000000000000000000000000000000000000;
				6'd56 : Enable_Registers <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
				6'd57 : Enable_Registers <= 64'b0000001000000000000000000000000000000000000000000000000000000000;
				6'd58 : Enable_Registers <= 64'b0000010000000000000000000000000000000000000000000000000000000000;
				6'd59 : Enable_Registers <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
				6'd60 : Enable_Registers <= 64'b0001000000000000000000000000000000000000000000000000000000000000;
				6'd61 : Enable_Registers <= 64'b0010000000000000000000000000000000000000000000000000000000000000;
				6'd62 : Enable_Registers <= 64'b0100000000000000000000000000000000000000000000000000000000000000;
				6'd63 : Enable_Registers <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_1024
	reg [4:0] Q_counter;
	reg [31:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset_TX_RX_Block | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset_TX_RX_Block | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				5'd0  : Enable_Registers <= 32'b00000000000000000000000000000001;
				5'd1  : Enable_Registers <= 32'b00000000000000000000000000000010;
				5'd2  : Enable_Registers <= 32'b00000000000000000000000000000100;
				5'd3  : Enable_Registers <= 32'b00000000000000000000000000001000;
				5'd4  : Enable_Registers <= 32'b00000000000000000000000000010000;
				5'd5  : Enable_Registers <= 32'b00000000000000000000000000100000;
				5'd6  : Enable_Registers <= 32'b00000000000000000000000001000000;
				5'd7  : Enable_Registers <= 32'b00000000000000000000000010000000;
				5'd8  : Enable_Registers <= 32'b00000000000000000000000100000000;
				5'd9  : Enable_Registers <= 32'b00000000000000000000001000000000;
				5'd10 : Enable_Registers <= 32'b00000000000000000000010000000000;
				5'd11 : Enable_Registers <= 32'b00000000000000000000100000000000;
				5'd12 : Enable_Registers <= 32'b00000000000000000001000000000000;
				5'd13 : Enable_Registers <= 32'b00000000000000000010000000000000;
				5'd14 : Enable_Registers <= 32'b00000000000000000100000000000000;
				5'd15 : Enable_Registers <= 32'b00000000000000001000000000000000;	
				5'd16 : Enable_Registers <= 32'b00000000000000010000000000000000;
				5'd17 : Enable_Registers <= 32'b00000000000000100000000000000000;
				5'd18 : Enable_Registers <= 32'b00000000000001000000000000000000;
				5'd19 : Enable_Registers <= 32'b00000000000010000000000000000000;
				5'd20 : Enable_Registers <= 32'b00000000000100000000000000000000;
				5'd21 : Enable_Registers <= 32'b00000000001000000000000000000000;
				5'd22 : Enable_Registers <= 32'b00000000010000000000000000000000;
				5'd23 : Enable_Registers <= 32'b00000000100000000000000000000000;
				5'd24 : Enable_Registers <= 32'b00000001000000000000000000000000;
				5'd25 : Enable_Registers <= 32'b00000010000000000000000000000000;
				5'd26 : Enable_Registers <= 32'b00000100000000000000000000000000;
				5'd27 : Enable_Registers <= 32'b00001000000000000000000000000000;
				5'd28 : Enable_Registers <= 32'b00010000000000000000000000000000;
				5'd29 : Enable_Registers <= 32'b00100000000000000000000000000000;
				5'd30 : Enable_Registers <= 32'b01000000000000000000000000000000;
				5'd31 : Enable_Registers <= 32'b10000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_512
	reg [3:0] Q_counter;
	reg [15:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				4'd0  : Enable_Registers <= 16'b0000000000000001;
				4'd1  : Enable_Registers <= 16'b0000000000000010;
				4'd2  : Enable_Registers <= 16'b0000000000000100;
				4'd3  : Enable_Registers <= 16'b0000000000001000;
				4'd4  : Enable_Registers <= 16'b0000000000010000;
				4'd5  : Enable_Registers <= 16'b0000000000100000;
				4'd6  : Enable_Registers <= 16'b0000000001000000;
				4'd7  : Enable_Registers <= 16'b0000000010000000;
				4'd8  : Enable_Registers <= 16'b0000000100000000;
				4'd9  : Enable_Registers <= 16'b0000001000000000;
				4'd10 : Enable_Registers <= 16'b0000010000000000;
				4'd11 : Enable_Registers <= 16'b0000100000000000;
				4'd12 : Enable_Registers <= 16'b0001000000000000;
				4'd13 : Enable_Registers <= 16'b0010000000000000;
				4'd14 : Enable_Registers <= 16'b0100000000000000;
				4'd15 : Enable_Registers <= 16'b1000000000000000;	
			endcase
`elsif PACKET_SIZE_256
	reg [2:0] Q_counter;
	reg [7:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter | reset_file_register)
				3'd0  : Enable_Registers <= 8'b00000001;
				3'd1  : Enable_Registers <= 8'b00000010;
				3'd2  : Enable_Registers <= 8'b00000100;
				3'd3  : Enable_Registers <= 8'b00001000;
				3'd4  : Enable_Registers <= 8'b00010000;
				3'd5  : Enable_Registers <= 8'b00100000;
				3'd6  : Enable_Registers <= 8'b01000000;
				3'd7  : Enable_Registers <= 8'b10000000;
			endcase
`elsif PACKET_SIZE_128
	reg [1:0] Q_counter;
	reg [3:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (reset | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (reset | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				2'd0  : Enable_Registers <= 4'b0001;
				2'd1  : Enable_Registers <= 4'b0010;
				2'd2  : Enable_Registers <= 4'b0100;
				2'd3  : Enable_Registers <= 4'b1000;
			endcase
`else
	// Statements
`endif

    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Máquina de estados finita
    // Se encarga del control de la ejecución de las acciones de este bloque.
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    

// ******************************************************  FSM *************************************************
	
	// Registro de estado
	always @(posedge user_clk) begin
	    if(reset_TX_RX_Block)
	        State<=S0;
	    else
	        State<=NextState;
	end
	
	// Lógica combinacional de estado siguiente
	always @* begin
	    case(State)
	            S0: begin  
                    NextState <= S1;
				end
				S1: begin // Wait for tlast               // Reset output register
                    if (m_axi_rx_tlast_reg) NextState <= S2;
            	    else NextState <= S1;
				end
				S2: begin // Wait for one clock cycle, for writing the last register in the register bank
                    NextState <= S3;
				end
				S3: begin // Load output register and reset all the register file and counter
					NextState <= S4;
                end	
				S4: begin // Wait if fifo is full and  Write wr_en flag is full is not asserted  
					if (full_reg) NextState <= S4;
            	    else NextState <= S1;
                end	
				default: begin 
					NextState <= S0;
                end				
		endcase
	end
                    	
	
	// Lógica combinacional de salida ************************************	
	always @* begin
	    case(State)
	           S0: begin  
                    reset_output_register <= 1'b1;
					wr_en_reg <= 1'b0;
					reset_file_register <= 1'b1;
					enable_output_register <= 1'b0;
				end
				S1: begin // Wait for tlast
                    reset_output_register <= 1'b1;
					wr_en_reg <= 1'b0;
					reset_file_register <= 1'b0;
					enable_output_register <= 1'b0;
				end
				S2: begin // Wait for the last write in the file register
					reset_output_register <= 1'b0;
					wr_en_reg <= 1'b0;
					reset_file_register <= 1'b0;
					enable_output_register <= 1'b0;
				end
				S3: begin // Load output register and reset all the register file and counter
					reset_output_register <= 1'b0;
					wr_en_reg <= 1'b0;
					reset_file_register <= 1'b1;
					enable_output_register <= 1'b1;
            end	
				S4: begin // Wait if fifo is full and  Write wr_en flag is full is not asserted  
					reset_output_register <= 1'b0;
					if (full_reg) wr_en_reg <= 1'b0;
            	    else wr_en_reg <= 1'b1;
					reset_file_register <= 1'b0;
					enable_output_register <= 1'b0;
            end	
				default: begin 
					reset_output_register <= 1'b1;
					wr_en_reg <= 1'b0;
					reset_file_register <= 1'b1;
					enable_output_register <= 1'b0;
            end				
		endcase
	end
	
	
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Memoria ROM
    // Se encarga de sustituir el secuenciador de paquetes por el BS_ID, para ello
    // toma como entrada el RX_UID (identificador global del nodo receptor) y genera
    // el identificador de BUS BS_ID
    // Se utiliza un parámetro definido como DATAFILE, el cual puede suponer valores válidos 
    // desde el 1 al 9. Esto sirve, ya que el DATAFILE varía en función de la FPGA donde
    // se encuentre.
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
    
    
	// ******************************************************  ROM Memory ******************************************
	
	ROM #(.DATAFILE(DATAFILE)) ROM_BS_UID(user_clk, din_reg[(PACKET_SIZE_BITS-1-32-8):(PACKET_SIZE_BITS-1-32-7-8)] , BS_ID);
	
	///////////////////////////////////////////////////////////////////////////////////////////////////
    // Registro de salida del paquete
    // Observe que este registro reemplaza el secuenciador de paquetes, por el 
    // BS_ID generado en la memoria ROM
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    
	register #(.WIDTH(PACKET_SIZE_BITS)) Parallel_Output_Register (
		.clk(user_clk), 
		.reset(reset_TX_RX_Block | reset_output_register), 
		.enable(enable_output_register), 
		.Din( {BS_ID, din_reg[PACKET_SIZE_BITS-1-8:0]} ), 
		.Dout(din)
	);
	
	
	// **************************************** Error handler
	
   ///////////////////////////////////////////////////////////////////////////////////////////////////
    // Contador de verificación de secuencia de paquete
    // Es un contador usado para verificación. El transmisor se encarga de colocar un
    // secuenciador de paquete, el cual se reemplaza en lugar del BS_ID, por su
    // parte el receptor, genera igualmente un secuenciador, pero para comparar
    // los datos con el secuenciador recibido, si estos difieren, significa que 
    // se rompió la secuencia de los paquetes y por ende, un error ocurrió.
    ///////////////////////////////////////////////////////////////////////////////////////////////////
    	
   
   always @(posedge user_clk)
      if (reset_TX_RX_Block)
         Q_seq_counter <= 0;
      else if (enable_output_register)
         Q_seq_counter <= Q_seq_counter + 1'b1;
	

   always @(posedge user_clk)
		if (reset_TX_RX_Block) begin
			Error <= 1'b0;
		end else if (Enable_Registers[1]) begin
			if (Q_seq_counter == din_reg[PACKET_SIZE_BITS-1:PACKET_SIZE_BITS-8])
				Error <= 1'b0;
			else
				Error <= 1'b1;
	   end

endmodule


module register #(parameter WIDTH = 32) (clk, reset, enable, Din, Dout);
    
    input clk, reset, enable;
    input [WIDTH-1:0] Din;
    output reg [WIDTH-1:0] Dout;
    
    always @(posedge clk) begin
        if (reset)
            Dout <= 0;
        else if (enable)
            Dout <= Din;
    end
    
endmodule

module ROM  #(parameter DATAFILE = 1) (CLK, Address, Output);
	
	localparam ROM_WIDTH = 8;
    localparam ROM_ADDR_BITS = 8;
	
	
	input CLK;
	input [ROM_ADDR_BITS-1:0] Address; // TX_UID 
	output reg [ROM_WIDTH-1:0] Output;  // BS_ID

   

    generate
        if (DATAFILE == 0) begin          // Esta memoria se usa en el ChannelTester_tb, Es un caso donde el Zynq está en el nodo 1.   
            always @(posedge CLK) 
                case (Address)
                    8'h00: Output <= 8'h01;
                    8'h01: Output <= 8'h01;
                    8'h02: Output <= 8'h01;
                    8'h03: Output <= 8'h01;
                    8'h04: Output <= 8'h01;
                    8'h05: Output <= 8'h01;
                    8'h06: Output <= 8'h01;
                    8'h07: Output <= 8'h01;
                    8'h08: Output <= 8'h01;
                    8'h09: Output <= 8'h01;
                    8'h0A: Output <= 8'h01;
                    8'h0B: Output <= 8'h01;
                    8'h0C: Output <= 8'h01;
                    8'h0D: Output <= 8'h01;
                    8'h0E: Output <= 8'h01;
                    8'h0F: Output <= 8'h01;
                    8'h10: Output <= 8'h01;
                    8'h11: Output <= 8'h01;
                    8'h12: Output <= 8'h01;
                    8'h13: Output <= 8'h01;
                    8'h14: Output <= 8'h01;
                    default: Output <= 8'hFF;
                endcase 
        end else if (DATAFILE == 1) begin    // Esta memoria se usa en el script_TO_Create_Vivado_Project, Es un caso donde el Zynq está en el nodo 2.   
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h02;
                    8'h01: Output <= 8'h02;
                    8'h02: Output <= 8'h02;
                    8'h03: Output <= 8'h02;
                    8'h04: Output <= 8'h02;
                    8'h05: Output <= 8'h02;
                    8'h06: Output <= 8'h02;
                    8'h07: Output <= 8'h02;
                    8'h08: Output <= 8'h02;
                    8'h09: Output <= 8'h02;
                    8'h0A: Output <= 8'h02;
                    8'h0B: Output <= 8'h02;
                    8'h0C: Output <= 8'h02;
                    8'h0D: Output <= 8'h02;
                    8'h0E: Output <= 8'h02;
                    8'h0F: Output <= 8'h02;
                    8'h10: Output <= 8'h02;
                    8'h11: Output <= 8'h02;
                    8'h12: Output <= 8'h02;
                    8'h13: Output <= 8'h02;
                    8'h14: Output <= 8'h02;
                    default: Output <= 8'hFF;
                endcase  
        end else if (DATAFILE == 2) begin    // Esta memoria se usa en el Testbench1, Es un caso donde el Zynq está en el nodo 4.
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h04;
                    8'h01: Output <= 8'h04;
                    8'h02: Output <= 8'h04;
                    8'h03: Output <= 8'h04;
                    8'h04: Output <= 8'h04;
                    8'h05: Output <= 8'h04;
                    8'h06: Output <= 8'h04;
                    8'h07: Output <= 8'h04;
                    8'h08: Output <= 8'h04;
                    8'h09: Output <= 8'h04;
                    8'h0A: Output <= 8'h04;
                    8'h0B: Output <= 8'h04;
                    8'h0C: Output <= 8'h04;
                    8'h0D: Output <= 8'h04;
                    8'h0E: Output <= 8'h04;
                    8'h0F: Output <= 8'h04;
                    8'h10: Output <= 8'h04;
                    8'h11: Output <= 8'h04;
                    8'h12: Output <= 8'h04;
                    8'h13: Output <= 8'h04;
                    8'h14: Output <= 8'h04;
                    default: Output <= 8'h04;
                endcase   
        end else if (DATAFILE == 3) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase  
        end else if (DATAFILE == 4) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase   
        end else if (DATAFILE == 5) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase   
        end else if (DATAFILE == 6) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase   
        end else if (DATAFILE == 7) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase  
        end else if (DATAFILE == 8) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase    
        end else if (DATAFILE == 9) begin    
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase    
        end else begin
            always @(posedge CLK)
                case (Address)
                    8'h00: Output <= 8'h00;
                    8'h01: Output <= 8'h00;
                    8'h02: Output <= 8'h00;
                    8'h03: Output <= 8'h00;
                    8'h04: Output <= 8'h00;
                    8'h05: Output <= 8'h00;
                    8'h06: Output <= 8'h00;
                    8'h07: Output <= 8'h00;
                    8'h08: Output <= 8'h00;
                    8'h09: Output <= 8'h00;
                    8'h0A: Output <= 8'h00;
                    8'h0B: Output <= 8'h00;
                    8'h0C: Output <= 8'h00;
                    8'h0D: Output <= 8'h00;
                    8'h0E: Output <= 8'h00;
                    8'h0F: Output <= 8'h00;
                    8'h10: Output <= 8'h00;
                    8'h11: Output <= 8'h00;
                    8'h12: Output <= 8'h00;
                    8'h13: Output <= 8'h00;
                    8'h14: Output <= 8'h00;
                    default: Output <= 8'h00;
                endcase   
        end
    endgenerate

  
        
endmodule

/*
module ROM  #(parameter DATAFILE = 1) (CLK, Address, Output);
	
	localparam ROM_WIDTH = 8;
    localparam ROM_ADDR_BITS = 8;
	
	
	input CLK;
	input [ROM_ADDR_BITS-1:0] Address; // RX_UID 
	output reg [ROM_WIDTH-1:0] Output;  // BS_ID

    (* rom_style="{distributed | block}" *)
    reg [ROM_WIDTH-1:0] ROM1 [(2**ROM_ADDR_BITS)-1:0];
    

    generate
        if (DATAFILE == 1) begin       
             initial
                $readmemh("Memory_Content_1.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 2) begin    
            initial
                $readmemh("Memory_Content_2.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 3) begin    
            initial
                $readmemh("Memory_Content_3.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 4) begin    
            initial
                $readmemh("Memory_Content_4.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 5) begin    
            initial
                $readmemh("Memory_Content_5.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 6) begin    
            initial
                $readmemh("Memory_Content_6.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 7) begin    
            initial
                $readmemh("Memory_Content_7.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 8) begin    
            initial
                $readmemh("Memory_Content_8.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else if (DATAFILE == 9) begin    
            initial
                $readmemh("Memory_Content_9.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end else begin
            initial
                $readmemh("Memory_Content_10.txt", ROM1, 0, (2**ROM_ADDR_BITS)-1);    
        end
    endgenerate

    always @(posedge CLK)
            Output <= ROM1[Address];
        
        
endmodule

*/
