`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/21/2021 02:19:29 AM
// Design Name: 
// Module Name: fifo_to_Aurora_One_lane_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fifo_to_Aurora_One_lane_tb;
    
    parameter PACKET_SIZE_BITS = 256; 
    //parameter PACKET_SIZE_BITS = 512; 
    //parameter PACKET_SIZE_BITS = 1024; 
    
    parameter NUMBER_OF_LANES = 1; 
    parameter ID_TARGET_FPGA = 8'h00;
    parameter n = 32*NUMBER_OF_LANES; 
    
    reg  user_clk, reset_TX_RX_Block;
    reg empty, s_axi_tx_tready;
    wire rd_en, s_axi_tx_tlast, s_axi_tx_tvalid; 
    
    reg [PACKET_SIZE_BITS-1: 0] dout;
    wire [n-1: 0] s_axi_tx_tdata;
    
    
    fifo_to_Aurora #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS), .NUMBER_OF_LANES(NUMBER_OF_LANES), .ID_TARGET_FPGA(ID_TARGET_FPGA)) uut(
    .user_clk(user_clk), 
    .reset_TX_RX_Block(reset_TX_RX_Block), 
    .empty(empty), 
    .rd_en(rd_en), 
    .dout(dout), 
    .s_axi_tx_tdata(s_axi_tx_tdata), 
    .s_axi_tx_tlast(s_axi_tx_tlast),
    .s_axi_tx_tready(s_axi_tx_tready), 
    .s_axi_tx_tvalid(s_axi_tx_tvalid)
    );
    
    initial begin
        user_clk = 0;
        reset_TX_RX_Block = 1;
        empty = 1;
        s_axi_tx_tready = 0;
        
        /* Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 1024 bits
        
        dout = 1024'h00000001_01000078_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E; 
        
        #40 empty = 0;
        s_axi_tx_tready = 1;
        
        #80 reset_TX_RX_Block = 0;
        
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 1024'h00010001_01000078_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        
        #32 empty = 0; 
        #32 empty = 1;
        #640 empty = 0; 
        #32 empty = 1;
        #640 empty = 0; 
        #32 empty = 1; 
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000078_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000074_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000070_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100006C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000068_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000064_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000060_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100005C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000058_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000054_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000050_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100004C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000048_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000044_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000040_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100003C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000038_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000034_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000030_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100002C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000028_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000024_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000020_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100001C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000018_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000014_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000010_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_0100000C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000008_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000004_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
        #640 empty = 0; 
       
        #640 s_axi_tx_tready = 0; 
        
        dout = 1024'h00010001_01000078_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D_0000001E;  
    
        #640 s_axi_tx_tready = 1; 
                                
        #2000 reset_TX_RX_Block = 1'b1;
        #80 reset_TX_RX_Block = 1'b0;
    
        // */
        
        /* Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 512 bits
        
        dout = 512'h00000001_01000038_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E; 
        
        
        #16 empty = 0;
        s_axi_tx_tready = 1; 
        
        #80 reset_TX_RX_Block = 0;
        
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 512'h00010001_01000038_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;  
        
        #32 empty = 0; 
        #32 empty = 1;
        #320 empty = 0; 
        #32 empty = 1;
        #320 empty = 0; 
        #32 empty = 1; 
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000034_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;  
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000030_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_0100002C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000028_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000024_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000020_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_0100001C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000018_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000014_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;  
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000010_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_0100000C_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000008_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000004_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E;   
        #320 empty = 0;         
        #320 s_axi_tx_tready = 0; 
        
        dout = 512'h00010001_01000038_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E; 
        #320 s_axi_tx_tready = 1;
        
        #320 dout = 512'h00010001_01000038_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E; 
        
        #1200 reset_TX_RX_Block = 1'b1;
        #80 reset_TX_RX_Block = 1'b0;
        
        // */
       
        
        // Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 256 bits
        
        
        dout = 256'h00000001_01000018_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #16 empty = 0;
        s_axi_tx_tready = 1; 
        
        
        #80 reset_TX_RX_Block = 0;
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 256'h00010001_01000018_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #32 empty = 0; 
        #32 empty = 1;
        #160 empty = 0; 
        #32 empty = 1;
        #160 empty = 0; 
        #32 empty = 1; 
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000014_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000010_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_0100000C_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000008_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000004_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        #160 empty = 0; 
         
        #160 s_axi_tx_tready = 0; 
        
        dout = 256'h00010001_01000018_00000001_00000002_00000003_00000004_00000005_00000006; 
    
        #160 s_axi_tx_tready = 1; 
        
        
        #200 dout = 256'h00010001_01000018_00000001_00000002_00000003_00000004_00000005_00000006; 
        
        
        #800 reset_TX_RX_Block = 1'b1;
        #80 reset_TX_RX_Block = 1'b0;
        
        
        // */
        
    end
    
    initial forever #4 user_clk = ~user_clk;


endmodule