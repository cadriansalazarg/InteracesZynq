`timescale 1ns / 1ps

`define PACKET_SIZE_256
//`define PACKET_SIZE_512
//`define PACKET_SIZE_1024

`ifdef PACKET_SIZE_256

    module FIFO_to_Custom_IP_tb;
        
        parameter PACKET_SIZE_BITS = 256;
        
        reg [PACKET_SIZE_BITS-1:0] dout;
        reg empty;
        wire rd_en;
            
        wire [7:0] in_fifo_V_BS_ID_dout;
        wire in_fifo_V_BS_ID_empty_n;
        reg in_fifo_V_BS_ID_read;
            
        wire [7:0] in_fifo_V_FPGA_ID_dout;
        wire in_fifo_V_FPGA_ID_empty_n;
            
        wire [15:0] in_fifo_V_PCKG_ID_dout;
        wire in_fifo_V_PCKG_ID_empty_n;
            
        wire [7:0] in_fifo_V_TX_UID_dout;
        wire in_fifo_V_TX_UID_empty_n;
            
        wire [7:0] in_fifo_V_RX_UID_dout;
        wire in_fifo_V_RX_UID_empty_n;
            
        wire [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        wire in_fifo_V_VALID_PACKET_BYTES_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_0_dout;
        wire in_fifo_V_MESSAGE_0_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_1_dout;
        wire in_fifo_V_MESSAGE_1_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_2_dout;
        wire in_fifo_V_MESSAGE_2_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_3_dout;
        wire in_fifo_V_MESSAGE_3_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_4_dout;
        wire in_fifo_V_MESSAGE_4_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_5_dout;
        wire in_fifo_V_MESSAGE_5_empty_n;
        
        FIFO_to_Custom_IP #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut (
            .rd_en(rd_en), 
            .dout(dout), 
            .empty(empty), 
            .in_fifo_V_BS_ID_dout(in_fifo_V_BS_ID_dout), 
            .in_fifo_V_BS_ID_empty_n(in_fifo_V_BS_ID_empty_n), 
            .in_fifo_V_BS_ID_read(in_fifo_V_BS_ID_read),
            .in_fifo_V_FPGA_ID_dout(in_fifo_V_FPGA_ID_dout), 
            .in_fifo_V_FPGA_ID_empty_n(in_fifo_V_FPGA_ID_empty_n),
            .in_fifo_V_PCKG_ID_dout(in_fifo_V_PCKG_ID_dout), 
            .in_fifo_V_PCKG_ID_empty_n(in_fifo_V_PCKG_ID_empty_n),
            .in_fifo_V_TX_UID_dout(in_fifo_V_TX_UID_dout), 
            .in_fifo_V_TX_UID_empty_n(in_fifo_V_TX_UID_empty_n),
            .in_fifo_V_RX_UID_dout(in_fifo_V_RX_UID_dout), 
            .in_fifo_V_RX_UID_empty_n(in_fifo_V_RX_UID_empty_n),
            .in_fifo_V_VALID_PACKET_BYTES_dout(in_fifo_V_VALID_PACKET_BYTES_dout), 
            .in_fifo_V_VALID_PACKET_BYTES_empty_n(in_fifo_V_VALID_PACKET_BYTES_empty_n),
            .in_fifo_V_MESSAGE_0_dout(in_fifo_V_MESSAGE_0_dout), 
            .in_fifo_V_MESSAGE_0_empty_n(in_fifo_V_MESSAGE_0_empty_n),
            .in_fifo_V_MESSAGE_1_dout(in_fifo_V_MESSAGE_1_dout), 
            .in_fifo_V_MESSAGE_1_empty_n(in_fifo_V_MESSAGE_1_empty_n),
            .in_fifo_V_MESSAGE_2_dout(in_fifo_V_MESSAGE_2_dout), 
            .in_fifo_V_MESSAGE_2_empty_n(in_fifo_V_MESSAGE_2_empty_n),
            .in_fifo_V_MESSAGE_3_dout(in_fifo_V_MESSAGE_3_dout), 
            .in_fifo_V_MESSAGE_3_empty_n(in_fifo_V_MESSAGE_3_empty_n),
            .in_fifo_V_MESSAGE_4_dout(in_fifo_V_MESSAGE_4_dout), 
            .in_fifo_V_MESSAGE_4_empty_n(in_fifo_V_MESSAGE_4_empty_n),
            .in_fifo_V_MESSAGE_5_dout(in_fifo_V_MESSAGE_5_dout), 
            .in_fifo_V_MESSAGE_5_empty_n(in_fifo_V_MESSAGE_5_empty_n)
        );
        
        initial begin
           
            dout = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            
            #400;
            dout = 256'h01234567_89ABCD0EF_00000000_00000001_00000002_00000003_00000004_00000005;
            
            #200;
            in_fifo_V_BS_ID_read = 1;
            
            #200;
            empty = 1;
            
            #20;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            dout = 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
            
            #400;
            empty = 1;
            in_fifo_V_BS_ID_read = 1;
            dout = 256'h01234567_89ABCD0EF_00000000_00000001_00000002_00000003_00000004_00000005;
    
            #400;
            dout = 256'hFFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF;
        end
    
    endmodule
    
`elsif PACKET_SIZE_512

    module FIFO_to_Custom_IP_tb;
        
        parameter PACKET_SIZE_BITS = 512;
        
        reg [PACKET_SIZE_BITS-1:0] dout;
        reg empty;
        wire rd_en;
            
        wire [7:0] in_fifo_V_BS_ID_dout;
        wire in_fifo_V_BS_ID_empty_n;
        reg in_fifo_V_BS_ID_read;
            
        wire [7:0] in_fifo_V_FPGA_ID_dout;
        wire in_fifo_V_FPGA_ID_empty_n;
            
        wire [15:0] in_fifo_V_PCKG_ID_dout;
        wire in_fifo_V_PCKG_ID_empty_n;
            
        wire [7:0] in_fifo_V_TX_UID_dout;
        wire in_fifo_V_TX_UID_empty_n;
            
        wire [7:0] in_fifo_V_RX_UID_dout;
        wire in_fifo_V_RX_UID_empty_n;
            
        wire [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        wire in_fifo_V_VALID_PACKET_BYTES_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_0_dout;
        wire in_fifo_V_MESSAGE_0_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_1_dout;
        wire in_fifo_V_MESSAGE_1_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_2_dout;
        wire in_fifo_V_MESSAGE_2_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_3_dout;
        wire in_fifo_V_MESSAGE_3_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_4_dout;
        wire in_fifo_V_MESSAGE_4_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_5_dout;
        wire in_fifo_V_MESSAGE_5_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_6_dout;
        wire in_fifo_V_MESSAGE_6_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_7_dout;
        wire in_fifo_V_MESSAGE_7_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_8_dout;
        wire in_fifo_V_MESSAGE_8_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_9_dout;
        wire in_fifo_V_MESSAGE_9_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_10_dout;
        wire in_fifo_V_MESSAGE_10_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_11_dout;
        wire in_fifo_V_MESSAGE_11_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_12_dout;
        wire in_fifo_V_MESSAGE_12_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_13_dout;
        wire in_fifo_V_MESSAGE_13_empty_n;
        
        FIFO_to_Custom_IP #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut (
            .rd_en(rd_en), 
            .dout(dout), 
            .empty(empty), 
            .in_fifo_V_BS_ID_dout(in_fifo_V_BS_ID_dout), 
            .in_fifo_V_BS_ID_empty_n(in_fifo_V_BS_ID_empty_n), 
            .in_fifo_V_BS_ID_read(in_fifo_V_BS_ID_read),
            .in_fifo_V_FPGA_ID_dout(in_fifo_V_FPGA_ID_dout), 
            .in_fifo_V_FPGA_ID_empty_n(in_fifo_V_FPGA_ID_empty_n),
            .in_fifo_V_PCKG_ID_dout(in_fifo_V_PCKG_ID_dout), 
            .in_fifo_V_PCKG_ID_empty_n(in_fifo_V_PCKG_ID_empty_n),
            .in_fifo_V_TX_UID_dout(in_fifo_V_TX_UID_dout), 
            .in_fifo_V_TX_UID_empty_n(in_fifo_V_TX_UID_empty_n),
            .in_fifo_V_RX_UID_dout(in_fifo_V_RX_UID_dout), 
            .in_fifo_V_RX_UID_empty_n(in_fifo_V_RX_UID_empty_n),
            .in_fifo_V_VALID_PACKET_BYTES_dout(in_fifo_V_VALID_PACKET_BYTES_dout), 
            .in_fifo_V_VALID_PACKET_BYTES_empty_n(in_fifo_V_VALID_PACKET_BYTES_empty_n),
            .in_fifo_V_MESSAGE_0_dout(in_fifo_V_MESSAGE_0_dout), 
            .in_fifo_V_MESSAGE_0_empty_n(in_fifo_V_MESSAGE_0_empty_n),
            .in_fifo_V_MESSAGE_1_dout(in_fifo_V_MESSAGE_1_dout), 
            .in_fifo_V_MESSAGE_1_empty_n(in_fifo_V_MESSAGE_1_empty_n),
            .in_fifo_V_MESSAGE_2_dout(in_fifo_V_MESSAGE_2_dout), 
            .in_fifo_V_MESSAGE_2_empty_n(in_fifo_V_MESSAGE_2_empty_n),
            .in_fifo_V_MESSAGE_3_dout(in_fifo_V_MESSAGE_3_dout), 
            .in_fifo_V_MESSAGE_3_empty_n(in_fifo_V_MESSAGE_3_empty_n),
            .in_fifo_V_MESSAGE_4_dout(in_fifo_V_MESSAGE_4_dout), 
            .in_fifo_V_MESSAGE_4_empty_n(in_fifo_V_MESSAGE_4_empty_n),
            .in_fifo_V_MESSAGE_5_dout(in_fifo_V_MESSAGE_5_dout), 
            .in_fifo_V_MESSAGE_5_empty_n(in_fifo_V_MESSAGE_5_empty_n),
            .in_fifo_V_MESSAGE_6_dout(in_fifo_V_MESSAGE_6_dout), 
            .in_fifo_V_MESSAGE_6_empty_n(in_fifo_V_MESSAGE_6_empty_n),
            .in_fifo_V_MESSAGE_7_dout(in_fifo_V_MESSAGE_7_dout), 
            .in_fifo_V_MESSAGE_7_empty_n(in_fifo_V_MESSAGE_7_empty_n),
            .in_fifo_V_MESSAGE_8_dout(in_fifo_V_MESSAGE_8_dout), 
            .in_fifo_V_MESSAGE_8_empty_n(in_fifo_V_MESSAGE_8_empty_n),
            .in_fifo_V_MESSAGE_9_dout(in_fifo_V_MESSAGE_9_dout), 
            .in_fifo_V_MESSAGE_9_empty_n(in_fifo_V_MESSAGE_9_empty_n),
            .in_fifo_V_MESSAGE_10_dout(in_fifo_V_MESSAGE_10_dout), 
            .in_fifo_V_MESSAGE_10_empty_n(in_fifo_V_MESSAGE_10_empty_n),
            .in_fifo_V_MESSAGE_11_dout(in_fifo_V_MESSAGE_11_dout), 
            .in_fifo_V_MESSAGE_11_empty_n(in_fifo_V_MESSAGE_11_empty_n),
            .in_fifo_V_MESSAGE_12_dout(in_fifo_V_MESSAGE_12_dout), 
            .in_fifo_V_MESSAGE_12_empty_n(in_fifo_V_MESSAGE_12_empty_n),
            .in_fifo_V_MESSAGE_13_dout(in_fifo_V_MESSAGE_13_dout), 
            .in_fifo_V_MESSAGE_13_empty_n(in_fifo_V_MESSAGE_13_empty_n)
        );
        
        initial begin
           
            dout = 512'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            
            #400;
            dout = 512'h01234567_89ABCD0EF_00000000_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D;
            
            #200;
            in_fifo_V_BS_ID_read = 1;
            
            #200;
            empty = 1;
            
            #20;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            
            #400;
            dout = 512'hFFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF;
               
        end
    
    endmodule

`elsif PACKET_SIZE_1024

    module FIFO_to_Custom_IP_tb;
        
        parameter PACKET_SIZE_BITS = 1024;
        
        reg [PACKET_SIZE_BITS-1:0] dout;
        reg empty;
        wire rd_en;
            
        wire [7:0] in_fifo_V_BS_ID_dout;
        wire in_fifo_V_BS_ID_empty_n;
        reg in_fifo_V_BS_ID_read;
            
        wire [7:0] in_fifo_V_FPGA_ID_dout;
        wire in_fifo_V_FPGA_ID_empty_n;
            
        wire [15:0] in_fifo_V_PCKG_ID_dout;
        wire in_fifo_V_PCKG_ID_empty_n;
            
        wire [7:0] in_fifo_V_TX_UID_dout;
        wire in_fifo_V_TX_UID_empty_n;
            
        wire [7:0] in_fifo_V_RX_UID_dout;
        wire in_fifo_V_RX_UID_empty_n;
            
        wire [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        wire in_fifo_V_VALID_PACKET_BYTES_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_0_dout;
        wire in_fifo_V_MESSAGE_0_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_1_dout;
        wire in_fifo_V_MESSAGE_1_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_2_dout;
        wire in_fifo_V_MESSAGE_2_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_3_dout;
        wire in_fifo_V_MESSAGE_3_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_4_dout;
        wire in_fifo_V_MESSAGE_4_empty_n;
            
        wire [31:0] in_fifo_V_MESSAGE_5_dout;
        wire in_fifo_V_MESSAGE_5_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_6_dout;
        wire in_fifo_V_MESSAGE_6_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_7_dout;
        wire in_fifo_V_MESSAGE_7_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_8_dout;
        wire in_fifo_V_MESSAGE_8_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_9_dout;
        wire in_fifo_V_MESSAGE_9_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_10_dout;
        wire in_fifo_V_MESSAGE_10_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_11_dout;
        wire in_fifo_V_MESSAGE_11_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_12_dout;
        wire in_fifo_V_MESSAGE_12_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_13_dout;
        wire in_fifo_V_MESSAGE_13_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_14_dout;
        wire in_fifo_V_MESSAGE_14_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_15_dout;
        wire in_fifo_V_MESSAGE_15_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_16_dout;
        wire in_fifo_V_MESSAGE_16_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_17_dout;
        wire in_fifo_V_MESSAGE_17_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_18_dout;
        wire in_fifo_V_MESSAGE_18_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_19_dout;
        wire in_fifo_V_MESSAGE_19_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_20_dout;
        wire in_fifo_V_MESSAGE_20_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_21_dout;
        wire in_fifo_V_MESSAGE_21_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_22_dout;
        wire in_fifo_V_MESSAGE_22_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_23_dout;
        wire in_fifo_V_MESSAGE_23_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_24_dout;
        wire in_fifo_V_MESSAGE_24_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_25_dout;
        wire in_fifo_V_MESSAGE_25_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_26_dout;
        wire in_fifo_V_MESSAGE_26_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_27_dout;
        wire in_fifo_V_MESSAGE_27_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_28_dout;
        wire in_fifo_V_MESSAGE_28_empty_n;
        
        wire [31:0] in_fifo_V_MESSAGE_29_dout;
        wire in_fifo_V_MESSAGE_29_empty_n;
        
        FIFO_to_Custom_IP #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut (
            .rd_en(rd_en), 
            .dout(dout), 
            .empty(empty), 
            .in_fifo_V_BS_ID_dout(in_fifo_V_BS_ID_dout), 
            .in_fifo_V_BS_ID_empty_n(in_fifo_V_BS_ID_empty_n), 
            .in_fifo_V_BS_ID_read(in_fifo_V_BS_ID_read),
            .in_fifo_V_FPGA_ID_dout(in_fifo_V_FPGA_ID_dout), 
            .in_fifo_V_FPGA_ID_empty_n(in_fifo_V_FPGA_ID_empty_n),
            .in_fifo_V_PCKG_ID_dout(in_fifo_V_PCKG_ID_dout), 
            .in_fifo_V_PCKG_ID_empty_n(in_fifo_V_PCKG_ID_empty_n),
            .in_fifo_V_TX_UID_dout(in_fifo_V_TX_UID_dout), 
            .in_fifo_V_TX_UID_empty_n(in_fifo_V_TX_UID_empty_n),
            .in_fifo_V_RX_UID_dout(in_fifo_V_RX_UID_dout), 
            .in_fifo_V_RX_UID_empty_n(in_fifo_V_RX_UID_empty_n),
            .in_fifo_V_VALID_PACKET_BYTES_dout(in_fifo_V_VALID_PACKET_BYTES_dout), 
            .in_fifo_V_VALID_PACKET_BYTES_empty_n(in_fifo_V_VALID_PACKET_BYTES_empty_n),
            .in_fifo_V_MESSAGE_0_dout(in_fifo_V_MESSAGE_0_dout), 
            .in_fifo_V_MESSAGE_0_empty_n(in_fifo_V_MESSAGE_0_empty_n),
            .in_fifo_V_MESSAGE_1_dout(in_fifo_V_MESSAGE_1_dout), 
            .in_fifo_V_MESSAGE_1_empty_n(in_fifo_V_MESSAGE_1_empty_n),
            .in_fifo_V_MESSAGE_2_dout(in_fifo_V_MESSAGE_2_dout), 
            .in_fifo_V_MESSAGE_2_empty_n(in_fifo_V_MESSAGE_2_empty_n),
            .in_fifo_V_MESSAGE_3_dout(in_fifo_V_MESSAGE_3_dout), 
            .in_fifo_V_MESSAGE_3_empty_n(in_fifo_V_MESSAGE_3_empty_n),
            .in_fifo_V_MESSAGE_4_dout(in_fifo_V_MESSAGE_4_dout), 
            .in_fifo_V_MESSAGE_4_empty_n(in_fifo_V_MESSAGE_4_empty_n),
            .in_fifo_V_MESSAGE_5_dout(in_fifo_V_MESSAGE_5_dout), 
            .in_fifo_V_MESSAGE_5_empty_n(in_fifo_V_MESSAGE_5_empty_n),
            .in_fifo_V_MESSAGE_6_dout(in_fifo_V_MESSAGE_6_dout), 
            .in_fifo_V_MESSAGE_6_empty_n(in_fifo_V_MESSAGE_6_empty_n),
            .in_fifo_V_MESSAGE_7_dout(in_fifo_V_MESSAGE_7_dout), 
            .in_fifo_V_MESSAGE_7_empty_n(in_fifo_V_MESSAGE_7_empty_n),
            .in_fifo_V_MESSAGE_8_dout(in_fifo_V_MESSAGE_8_dout), 
            .in_fifo_V_MESSAGE_8_empty_n(in_fifo_V_MESSAGE_8_empty_n),
            .in_fifo_V_MESSAGE_9_dout(in_fifo_V_MESSAGE_9_dout), 
            .in_fifo_V_MESSAGE_9_empty_n(in_fifo_V_MESSAGE_9_empty_n),
            .in_fifo_V_MESSAGE_10_dout(in_fifo_V_MESSAGE_10_dout), 
            .in_fifo_V_MESSAGE_10_empty_n(in_fifo_V_MESSAGE_10_empty_n),
            .in_fifo_V_MESSAGE_11_dout(in_fifo_V_MESSAGE_11_dout), 
            .in_fifo_V_MESSAGE_11_empty_n(in_fifo_V_MESSAGE_11_empty_n),
            .in_fifo_V_MESSAGE_12_dout(in_fifo_V_MESSAGE_12_dout), 
            .in_fifo_V_MESSAGE_12_empty_n(in_fifo_V_MESSAGE_12_empty_n),
            .in_fifo_V_MESSAGE_13_dout(in_fifo_V_MESSAGE_13_dout), 
            .in_fifo_V_MESSAGE_13_empty_n(in_fifo_V_MESSAGE_13_empty_n),
            .in_fifo_V_MESSAGE_14_dout(in_fifo_V_MESSAGE_14_dout), 
            .in_fifo_V_MESSAGE_14_empty_n(in_fifo_V_MESSAGE_14_empty_n),
            .in_fifo_V_MESSAGE_15_dout(in_fifo_V_MESSAGE_15_dout), 
            .in_fifo_V_MESSAGE_15_empty_n(in_fifo_V_MESSAGE_15_empty_n),
            .in_fifo_V_MESSAGE_16_dout(in_fifo_V_MESSAGE_16_dout), 
            .in_fifo_V_MESSAGE_16_empty_n(in_fifo_V_MESSAGE_16_empty_n),
            .in_fifo_V_MESSAGE_17_dout(in_fifo_V_MESSAGE_17_dout), 
            .in_fifo_V_MESSAGE_17_empty_n(in_fifo_V_MESSAGE_17_empty_n),
            .in_fifo_V_MESSAGE_18_dout(in_fifo_V_MESSAGE_18_dout), 
            .in_fifo_V_MESSAGE_18_empty_n(in_fifo_V_MESSAGE_18_empty_n),
            .in_fifo_V_MESSAGE_19_dout(in_fifo_V_MESSAGE_19_dout), 
            .in_fifo_V_MESSAGE_19_empty_n(in_fifo_V_MESSAGE_19_empty_n),
            .in_fifo_V_MESSAGE_20_dout(in_fifo_V_MESSAGE_20_dout), 
            .in_fifo_V_MESSAGE_20_empty_n(in_fifo_V_MESSAGE_20_empty_n),
            .in_fifo_V_MESSAGE_21_dout(in_fifo_V_MESSAGE_21_dout), 
            .in_fifo_V_MESSAGE_21_empty_n(in_fifo_V_MESSAGE_21_empty_n),
            .in_fifo_V_MESSAGE_22_dout(in_fifo_V_MESSAGE_22_dout), 
            .in_fifo_V_MESSAGE_22_empty_n(in_fifo_V_MESSAGE_22_empty_n),
            .in_fifo_V_MESSAGE_23_dout(in_fifo_V_MESSAGE_23_dout), 
            .in_fifo_V_MESSAGE_23_empty_n(in_fifo_V_MESSAGE_23_empty_n),
            .in_fifo_V_MESSAGE_24_dout(in_fifo_V_MESSAGE_24_dout), 
            .in_fifo_V_MESSAGE_24_empty_n(in_fifo_V_MESSAGE_24_empty_n),
            .in_fifo_V_MESSAGE_25_dout(in_fifo_V_MESSAGE_25_dout), 
            .in_fifo_V_MESSAGE_25_empty_n(in_fifo_V_MESSAGE_25_empty_n),
            .in_fifo_V_MESSAGE_26_dout(in_fifo_V_MESSAGE_26_dout), 
            .in_fifo_V_MESSAGE_26_empty_n(in_fifo_V_MESSAGE_26_empty_n),
            .in_fifo_V_MESSAGE_27_dout(in_fifo_V_MESSAGE_27_dout), 
            .in_fifo_V_MESSAGE_27_empty_n(in_fifo_V_MESSAGE_27_empty_n),
            .in_fifo_V_MESSAGE_28_dout(in_fifo_V_MESSAGE_28_dout), 
            .in_fifo_V_MESSAGE_28_empty_n(in_fifo_V_MESSAGE_28_empty_n),
            .in_fifo_V_MESSAGE_29_dout(in_fifo_V_MESSAGE_29_dout), 
            .in_fifo_V_MESSAGE_29_empty_n(in_fifo_V_MESSAGE_29_empty_n)
        );
        
        initial begin
           
            dout = 1024'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            
            #400;
            dout = 1024'h01234567_89ABCDEF_00000000_00000001_00000002_00000003_00000004_00000005_00000006_00000007_00000008_00000009_0000000A_0000000B_0000000C_0000000D_0000000E_0000000F_00000010_00000011_00000012_00000013_00000014_00000015_00000016_00000017_00000018_00000019_0000001A_0000001B_0000001C_0000001D;
            
            #200;
            in_fifo_V_BS_ID_read = 1;
            
            #200;
            empty = 1;
            
            #20;
            empty = 0;
            in_fifo_V_BS_ID_read = 0;
            
            #400;
            dout = 1024'hFFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF;
               
        end
    
    endmodule


`else
	// Statements
`endif 