`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/21/2021 03:27:57 AM
// Design Name: 
// Module Name: fifo_to_Aurora_Two_lanes_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fifo_to_Aurora_Two_lanes_tb;
    
    //parameter PACKET_SIZE_BITS = 256; 
    //parameter PACKET_SIZE_BITS = 512; 
    parameter PACKET_SIZE_BITS = 1024; 
    
    parameter NUMBER_OF_LANES = 2; 
    parameter ID_TARGET_FPGA = 8'h00;
    parameter n = 32*NUMBER_OF_LANES; 
    
    reg  user_clk, reset_TX_RX_Block;
    reg empty, s_axi_tx_tready;
    wire rd_en, s_axi_tx_tlast, s_axi_tx_tvalid; 
    
    reg [PACKET_SIZE_BITS-1: 0] dout;
    wire [n-1: 0] s_axi_tx_tdata;
    
    
    fifo_to_Aurora #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS), .NUMBER_OF_LANES(NUMBER_OF_LANES), .ID_TARGET_FPGA(ID_TARGET_FPGA)) uut(
    .user_clk(user_clk), 
    .reset_TX_RX_Block(reset_TX_RX_Block), 
    .empty(empty), 
    .rd_en(rd_en), 
    .dout(dout), 
    .s_axi_tx_tdata(s_axi_tx_tdata), 
    .s_axi_tx_tlast(s_axi_tx_tlast),
    .s_axi_tx_tready(s_axi_tx_tready), 
    .s_axi_tx_tvalid(s_axi_tx_tvalid)
    );
    
    initial begin
        user_clk = 0;
        reset_TX_RX_Block = 1;
        empty = 1;
        s_axi_tx_tready = 0;
        
        // Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 1024 bits
        
        dout = 1024'h00000001_01000078_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F; 
        
        #160 empty = 0;
        s_axi_tx_tready = 1;
        
        #80 reset_TX_RX_Block = 0;
        
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 1024'h00010001_01000078_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        
        #32 empty = 0; 
        #32 empty = 1;
        #640 empty = 0; 
        #32 empty = 1;
        #640 empty = 0; 
        #32 empty = 1; 
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000078_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000070_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000068__00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000060_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000058_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000050_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000048_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000040_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000038_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000030_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000028_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000020_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000018_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000010_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #32 empty = 1;
        
        dout = 1024'h00010001_01000008_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
        #640 empty = 0; 
        #640 s_axi_tx_tready = 0; 
        
        dout = 1024'h00010001_01000078_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F;
    
        #640 s_axi_tx_tready = 1; 
        
        #640 dout = 1024'h00010001_01000078_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007_00000000_00000008_00000000_00000009_00000000_0000000A_00000000_0000000B_00000000_0000000C_00000000_0000000D_00000000_0000000E_00000000_0000000F; 
        
        #400 reset_TX_RX_Block = 1;
        
        #80 reset_TX_RX_Block = 0;
    
        // */
        
        /* Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 512 bits
        
        dout = 512'h00000001_01000038_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007; 
        
        #160 empty = 0;
        s_axi_tx_tready = 1;
        
        #80 reset_TX_RX_Block = 0;

        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 512'h00010001_01000038_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        
        #32 empty = 0; 
        #32 empty = 1;
        #320 empty = 0; 
        #32 empty = 1;
        #320 empty = 0; 
        #32 empty = 1; 
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000030_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
        #32 empty = 1;
               
        dout = 512'h00010001_01000028_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000020_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000018_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
        #32 empty = 1;
                
        dout = 512'h00010001_01000010_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
        #32 empty = 1;
        
        dout = 512'h00010001_01000008_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        #320 empty = 0; 
                
        #320 s_axi_tx_tready = 0; 
        
        dout = 512'h00010001_01000038_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
    
        #320 s_axi_tx_tready = 1; 
        #32 s_axi_tx_tready = 0;
        
        #320 s_axi_tx_tready = 1;
        
        #320 dout = 512'h00010001_01000038_00000000_00000001_00000000_00000002_00000000_00000003_00000000_00000004_00000000_00000005_00000000_00000006_00000000_00000007;
        
        #400 reset_TX_RX_Block = 1;
        
        #80 reset_TX_RX_Block = 0;
        // */
       
        
        /* Descomentar esta línea para verificar el funcionamiento de la versión con tamaño de paquete de 256 bits
        
        dout = 256'h00000001_01000018_00000000_00000001_00000000_00000002_00000000_00000003; 
        
        #160 empty = 0;
        s_axi_tx_tready = 1;
        
        #80 reset_TX_RX_Block = 0;
        
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        #32 empty = 0; 
        #32 empty = 1; 
        
        dout = 256'h00010001_01000018_00000000_00000001_00000000_00000002_00000000_00000003; 
        
        #32 empty = 0; 
        #32 empty = 1;
        #160 empty = 0; 
        #32 empty = 1;
        #160 empty = 0; 
        #32 empty = 1; 
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000010_00000000_00000001_00000000_00000002_00000000_00000003; 
        
        #160 empty = 0; 
        #32 empty = 1;
        
        dout = 256'h00010001_01000008_00000000_00000001_00000000_00000002_00000000_00000003; 
        
        #160 empty = 0; 
        
        #160 s_axi_tx_tready = 0; 
        
        dout = 256'h00010001_01000018_00000000_00000001_00000000_00000002_00000000_00000003; 
    
        #160 s_axi_tx_tready = 1; 
        #32 s_axi_tx_tready = 0;
        
        #160 s_axi_tx_tready = 1;
        
        #200 dout = 256'h00010001_01000018_00000000_00000001_00000000_00000002_00000000_00000003; 
        
        #400 reset_TX_RX_Block = 1;
        
        #80 reset_TX_RX_Block = 0;
        
        // */
        
    end
    
    initial forever #4 user_clk = ~user_clk;


endmodule