`timescale 1ns / 1ps

`define PACKET_SIZE_256
//`define PACKET_SIZE_512
//`define PACKET_SIZE_1024

`ifdef PACKET_SIZE_256

    module Custom_IP_to_FIFO_tb;
        
        parameter PACKET_SIZE_BITS = 256;
        
        wire wr_en;
        wire full_n;
        wire [PACKET_SIZE_BITS-1:0] din;
            
            
        reg [7:0] out_fifo_V_BS_ID_din;
        reg out_fifo_V_BS_ID_write;
        reg full;
            
        reg [7:0] out_fifo_V_FPGA_ID_din;
        reg [15:0] out_fifo_V_PCKG_ID_din;
        reg [7:0] out_fifo_V_TX_UID_din;
        reg [7:0] out_fifo_V_RX_UID_din;
        reg [15:0] out_fifo_V_VALID_PACKET_BYTES_din;
            
        reg [31:0] out_fifo_V_MESSAGE_0_din;
        reg [31:0] out_fifo_V_MESSAGE_1_din;
        reg [31:0] out_fifo_V_MESSAGE_2_din;
        reg [31:0] out_fifo_V_MESSAGE_3_din;
        reg [31:0] out_fifo_V_MESSAGE_4_din;
        reg [31:0] out_fifo_V_MESSAGE_5_din; 
        
        Custom_IP_to_FIFO #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut(
            .wr_en(wr_en), 
            .din(din), 
            .full(full),
            .full_n(full_n),
            .out_fifo_V_BS_ID_din(out_fifo_V_BS_ID_din), 
            .out_fifo_V_BS_ID_write(out_fifo_V_BS_ID_write),
            .out_fifo_V_FPGA_ID_din(out_fifo_V_FPGA_ID_din),
            .out_fifo_V_PCKG_ID_din(out_fifo_V_PCKG_ID_din), 
            .out_fifo_V_TX_UID_din(out_fifo_V_TX_UID_din),
            .out_fifo_V_RX_UID_din(out_fifo_V_RX_UID_din), 
            .out_fifo_V_VALID_PACKET_BYTES_din(out_fifo_V_VALID_PACKET_BYTES_din),
            .out_fifo_V_MESSAGE_0_din(out_fifo_V_MESSAGE_0_din),
            .out_fifo_V_MESSAGE_1_din(out_fifo_V_MESSAGE_1_din), 
            .out_fifo_V_MESSAGE_2_din(out_fifo_V_MESSAGE_2_din), 
            .out_fifo_V_MESSAGE_3_din(out_fifo_V_MESSAGE_3_din), 
            .out_fifo_V_MESSAGE_4_din(out_fifo_V_MESSAGE_4_din), 
            .out_fifo_V_MESSAGE_5_din(out_fifo_V_MESSAGE_5_din) 
        );
        
        initial begin
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            full = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'hFF;
            out_fifo_V_BS_ID_write = 1;
            full = 1;
            
            out_fifo_V_FPGA_ID_din = 8'hFF;
            out_fifo_V_PCKG_ID_din = 16'hFFFF;
            out_fifo_V_TX_UID_din = 8'hFF;
            out_fifo_V_RX_UID_din = 8'hFF;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'hFFFE;
            
            out_fifo_V_MESSAGE_0_din = 32'hFFFFFFFD;
            out_fifo_V_MESSAGE_1_din = 32'hFFFFFFFC;
            out_fifo_V_MESSAGE_2_din = 32'hFFFFFFFB;
            out_fifo_V_MESSAGE_3_din = 32'hFFFFFFFA;
            out_fifo_V_MESSAGE_4_din = 32'hFFFFFFF9;
            out_fifo_V_MESSAGE_5_din = 32'hFFFFFFF8;
            
            #400;
            
            
            #200;
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0000;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000000;
            out_fifo_V_MESSAGE_1_din = 32'h00000000;
            out_fifo_V_MESSAGE_2_din = 32'h00000000;
            out_fifo_V_MESSAGE_3_din = 32'h00000000;
            out_fifo_V_MESSAGE_4_din = 32'h00000000;
            out_fifo_V_MESSAGE_5_din = 32'h00000000;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 1;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            
        end
        
    
    endmodule

`elsif PACKET_SIZE_512

    module Custom_IP_to_FIFO_tb;
        
        parameter PACKET_SIZE_BITS = 512;
        
        wire wr_en, full_n;
        wire [PACKET_SIZE_BITS-1:0] din;
            
            
        reg [7:0] out_fifo_V_BS_ID_din;
        reg out_fifo_V_BS_ID_write;
        reg full;
            
        reg [7:0] out_fifo_V_FPGA_ID_din;
        reg [15:0] out_fifo_V_PCKG_ID_din;
        reg [7:0] out_fifo_V_TX_UID_din;
        reg [7:0] out_fifo_V_RX_UID_din;
        reg [15:0] out_fifo_V_VALID_PACKET_BYTES_din;
            
        reg [31:0] out_fifo_V_MESSAGE_0_din;
        reg [31:0] out_fifo_V_MESSAGE_1_din;
        reg [31:0] out_fifo_V_MESSAGE_2_din;
        reg [31:0] out_fifo_V_MESSAGE_3_din;
        reg [31:0] out_fifo_V_MESSAGE_4_din;
        reg [31:0] out_fifo_V_MESSAGE_5_din; 
        reg [31:0] out_fifo_V_MESSAGE_6_din; 
        reg [31:0] out_fifo_V_MESSAGE_7_din; 
        reg [31:0] out_fifo_V_MESSAGE_8_din; 
        reg [31:0] out_fifo_V_MESSAGE_9_din; 
        reg [31:0] out_fifo_V_MESSAGE_10_din; 
        reg [31:0] out_fifo_V_MESSAGE_11_din; 
        reg [31:0] out_fifo_V_MESSAGE_12_din; 
        reg [31:0] out_fifo_V_MESSAGE_13_din; 
        
        Custom_IP_to_FIFO #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut(
            .wr_en(wr_en), 
            .din(din), 
            .full(full),
            .full_n(full_n),
            .out_fifo_V_BS_ID_din(out_fifo_V_BS_ID_din), 
            .out_fifo_V_BS_ID_write(out_fifo_V_BS_ID_write),
            .out_fifo_V_FPGA_ID_din(out_fifo_V_FPGA_ID_din),
            .out_fifo_V_PCKG_ID_din(out_fifo_V_PCKG_ID_din), 
            .out_fifo_V_TX_UID_din(out_fifo_V_TX_UID_din),
            .out_fifo_V_RX_UID_din(out_fifo_V_RX_UID_din), 
            .out_fifo_V_VALID_PACKET_BYTES_din(out_fifo_V_VALID_PACKET_BYTES_din),
            .out_fifo_V_MESSAGE_0_din(out_fifo_V_MESSAGE_0_din),
            .out_fifo_V_MESSAGE_1_din(out_fifo_V_MESSAGE_1_din), 
            .out_fifo_V_MESSAGE_2_din(out_fifo_V_MESSAGE_2_din), 
            .out_fifo_V_MESSAGE_3_din(out_fifo_V_MESSAGE_3_din), 
            .out_fifo_V_MESSAGE_4_din(out_fifo_V_MESSAGE_4_din), 
            .out_fifo_V_MESSAGE_5_din(out_fifo_V_MESSAGE_5_din),
            .out_fifo_V_MESSAGE_6_din(out_fifo_V_MESSAGE_6_din), 
            .out_fifo_V_MESSAGE_7_din(out_fifo_V_MESSAGE_7_din), 
            .out_fifo_V_MESSAGE_8_din(out_fifo_V_MESSAGE_8_din), 
            .out_fifo_V_MESSAGE_9_din(out_fifo_V_MESSAGE_9_din), 
            .out_fifo_V_MESSAGE_10_din(out_fifo_V_MESSAGE_10_din), 
            .out_fifo_V_MESSAGE_11_din(out_fifo_V_MESSAGE_11_din), 
            .out_fifo_V_MESSAGE_12_din(out_fifo_V_MESSAGE_12_din), 
            .out_fifo_V_MESSAGE_13_din(out_fifo_V_MESSAGE_13_din)             
        );
        
        initial begin
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            full = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            out_fifo_V_MESSAGE_6_din = 32'h00000008;
            out_fifo_V_MESSAGE_7_din = 32'h00000009;
            out_fifo_V_MESSAGE_8_din = 32'h0000000A;
            out_fifo_V_MESSAGE_9_din = 32'h0000000B;
            out_fifo_V_MESSAGE_10_din = 32'h0000000C;
            out_fifo_V_MESSAGE_11_din = 32'h0000000D;
            out_fifo_V_MESSAGE_12_din = 32'h0000000E;
            out_fifo_V_MESSAGE_13_din = 32'h0000000F;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'hFF;
            out_fifo_V_BS_ID_write = 1;
            full = 1;
            
            out_fifo_V_FPGA_ID_din = 8'hFF;
            out_fifo_V_PCKG_ID_din = 16'hFFFF;
            out_fifo_V_TX_UID_din = 8'hFF;
            out_fifo_V_RX_UID_din = 8'hFF;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'hFFFE;
            
            out_fifo_V_MESSAGE_0_din = 32'hFFFFFFFD;
            out_fifo_V_MESSAGE_1_din = 32'hFFFFFFFC;
            out_fifo_V_MESSAGE_2_din = 32'hFFFFFFFB;
            out_fifo_V_MESSAGE_3_din = 32'hFFFFFFFA;
            out_fifo_V_MESSAGE_4_din = 32'hFFFFFFF9;
            out_fifo_V_MESSAGE_5_din = 32'hFFFFFFF8;
            out_fifo_V_MESSAGE_6_din = 32'hFFFFFFF7;
            out_fifo_V_MESSAGE_7_din = 32'hFFFFFFF6;
            out_fifo_V_MESSAGE_8_din = 32'hFFFFFFF5;
            out_fifo_V_MESSAGE_9_din = 32'hFFFFFFF4;
            out_fifo_V_MESSAGE_10_din = 32'hFFFFFFF3;
            out_fifo_V_MESSAGE_11_din = 32'hFFFFFFF2;
            out_fifo_V_MESSAGE_12_din = 32'hFFFFFFF1;
            out_fifo_V_MESSAGE_13_din = 32'hFFFFFFF0;
            
            
            #200;
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0000;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000000;
            out_fifo_V_MESSAGE_1_din = 32'h00000000;
            out_fifo_V_MESSAGE_2_din = 32'h00000000;
            out_fifo_V_MESSAGE_3_din = 32'h00000000;
            out_fifo_V_MESSAGE_4_din = 32'h00000000;
            out_fifo_V_MESSAGE_5_din = 32'h00000000;
            out_fifo_V_MESSAGE_6_din = 32'h00000000;
            out_fifo_V_MESSAGE_7_din = 32'h00000000;
            out_fifo_V_MESSAGE_8_din = 32'h00000000;
            out_fifo_V_MESSAGE_9_din = 32'h00000000;
            out_fifo_V_MESSAGE_10_din = 32'h00000000;
            out_fifo_V_MESSAGE_11_din = 32'h00000000;
            out_fifo_V_MESSAGE_12_din = 32'h00000000;
            out_fifo_V_MESSAGE_13_din = 32'h00000000;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 1;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            out_fifo_V_MESSAGE_6_din = 32'h00000008;
            out_fifo_V_MESSAGE_7_din = 32'h00000009;
            out_fifo_V_MESSAGE_8_din = 32'h0000000A;
            out_fifo_V_MESSAGE_9_din = 32'h0000000B;
            out_fifo_V_MESSAGE_10_din = 32'h0000000C;
            out_fifo_V_MESSAGE_11_din = 32'h0000000D;
            out_fifo_V_MESSAGE_12_din = 32'h0000000E;
            out_fifo_V_MESSAGE_13_din = 32'h0000000F;
            
        end
            
    endmodule

`elsif PACKET_SIZE_1024 

    module Custom_IP_to_FIFO_tb;
        
        parameter PACKET_SIZE_BITS = 1024;
        
        wire wr_en, full_n;
        wire [PACKET_SIZE_BITS-1:0] din;
            
            
        reg [7:0] out_fifo_V_BS_ID_din;
        reg out_fifo_V_BS_ID_write;
        reg full;
            
        reg [7:0] out_fifo_V_FPGA_ID_din;
        reg [15:0] out_fifo_V_PCKG_ID_din;
        reg [7:0] out_fifo_V_TX_UID_din;
        reg [7:0] out_fifo_V_RX_UID_din;
        reg [15:0] out_fifo_V_VALID_PACKET_BYTES_din;
            
        reg [31:0] out_fifo_V_MESSAGE_0_din;
        reg [31:0] out_fifo_V_MESSAGE_1_din;
        reg [31:0] out_fifo_V_MESSAGE_2_din;
        reg [31:0] out_fifo_V_MESSAGE_3_din;
        reg [31:0] out_fifo_V_MESSAGE_4_din;
        reg [31:0] out_fifo_V_MESSAGE_5_din; 
        reg [31:0] out_fifo_V_MESSAGE_6_din; 
        reg [31:0] out_fifo_V_MESSAGE_7_din; 
        reg [31:0] out_fifo_V_MESSAGE_8_din; 
        reg [31:0] out_fifo_V_MESSAGE_9_din; 
        reg [31:0] out_fifo_V_MESSAGE_10_din; 
        reg [31:0] out_fifo_V_MESSAGE_11_din; 
        reg [31:0] out_fifo_V_MESSAGE_12_din; 
        reg [31:0] out_fifo_V_MESSAGE_13_din; 
        reg [31:0] out_fifo_V_MESSAGE_14_din;
        reg [31:0] out_fifo_V_MESSAGE_15_din;
        reg [31:0] out_fifo_V_MESSAGE_16_din;
        reg [31:0] out_fifo_V_MESSAGE_17_din;
        reg [31:0] out_fifo_V_MESSAGE_18_din;
        reg [31:0] out_fifo_V_MESSAGE_19_din;
        reg [31:0] out_fifo_V_MESSAGE_20_din;
        reg [31:0] out_fifo_V_MESSAGE_21_din;
        reg [31:0] out_fifo_V_MESSAGE_22_din;
        reg [31:0] out_fifo_V_MESSAGE_23_din;
        reg [31:0] out_fifo_V_MESSAGE_24_din;
        reg [31:0] out_fifo_V_MESSAGE_25_din;
        reg [31:0] out_fifo_V_MESSAGE_26_din;
        reg [31:0] out_fifo_V_MESSAGE_27_din;
        reg [31:0] out_fifo_V_MESSAGE_28_din;
        reg [31:0] out_fifo_V_MESSAGE_29_din;
        
        Custom_IP_to_FIFO #(.PACKET_SIZE_BITS(PACKET_SIZE_BITS)) uut(
            .wr_en(wr_en), 
            .din(din), 
            .full(full),
            .full_n(full_n),
            .out_fifo_V_BS_ID_din(out_fifo_V_BS_ID_din), 
            .out_fifo_V_BS_ID_write(out_fifo_V_BS_ID_write),
            .out_fifo_V_FPGA_ID_din(out_fifo_V_FPGA_ID_din),
            .out_fifo_V_PCKG_ID_din(out_fifo_V_PCKG_ID_din), 
            .out_fifo_V_TX_UID_din(out_fifo_V_TX_UID_din),
            .out_fifo_V_RX_UID_din(out_fifo_V_RX_UID_din), 
            .out_fifo_V_VALID_PACKET_BYTES_din(out_fifo_V_VALID_PACKET_BYTES_din),
            .out_fifo_V_MESSAGE_0_din(out_fifo_V_MESSAGE_0_din),
            .out_fifo_V_MESSAGE_1_din(out_fifo_V_MESSAGE_1_din), 
            .out_fifo_V_MESSAGE_2_din(out_fifo_V_MESSAGE_2_din), 
            .out_fifo_V_MESSAGE_3_din(out_fifo_V_MESSAGE_3_din), 
            .out_fifo_V_MESSAGE_4_din(out_fifo_V_MESSAGE_4_din), 
            .out_fifo_V_MESSAGE_5_din(out_fifo_V_MESSAGE_5_din),
            .out_fifo_V_MESSAGE_6_din(out_fifo_V_MESSAGE_6_din), 
            .out_fifo_V_MESSAGE_7_din(out_fifo_V_MESSAGE_7_din), 
            .out_fifo_V_MESSAGE_8_din(out_fifo_V_MESSAGE_8_din), 
            .out_fifo_V_MESSAGE_9_din(out_fifo_V_MESSAGE_9_din), 
            .out_fifo_V_MESSAGE_10_din(out_fifo_V_MESSAGE_10_din), 
            .out_fifo_V_MESSAGE_11_din(out_fifo_V_MESSAGE_11_din), 
            .out_fifo_V_MESSAGE_12_din(out_fifo_V_MESSAGE_12_din), 
            .out_fifo_V_MESSAGE_13_din(out_fifo_V_MESSAGE_13_din),  
            .out_fifo_V_MESSAGE_14_din(out_fifo_V_MESSAGE_14_din), 
            .out_fifo_V_MESSAGE_15_din(out_fifo_V_MESSAGE_15_din), 
            .out_fifo_V_MESSAGE_16_din(out_fifo_V_MESSAGE_16_din), 
            .out_fifo_V_MESSAGE_17_din(out_fifo_V_MESSAGE_17_din), 
            .out_fifo_V_MESSAGE_18_din(out_fifo_V_MESSAGE_18_din), 
            .out_fifo_V_MESSAGE_19_din(out_fifo_V_MESSAGE_19_din), 
            .out_fifo_V_MESSAGE_20_din(out_fifo_V_MESSAGE_20_din), 
            .out_fifo_V_MESSAGE_21_din(out_fifo_V_MESSAGE_21_din), 
            .out_fifo_V_MESSAGE_22_din(out_fifo_V_MESSAGE_22_din), 
            .out_fifo_V_MESSAGE_23_din(out_fifo_V_MESSAGE_23_din), 
            .out_fifo_V_MESSAGE_24_din(out_fifo_V_MESSAGE_24_din), 
            .out_fifo_V_MESSAGE_25_din(out_fifo_V_MESSAGE_25_din), 
            .out_fifo_V_MESSAGE_26_din(out_fifo_V_MESSAGE_26_din), 
            .out_fifo_V_MESSAGE_27_din(out_fifo_V_MESSAGE_27_din), 
            .out_fifo_V_MESSAGE_28_din(out_fifo_V_MESSAGE_28_din), 
            .out_fifo_V_MESSAGE_29_din(out_fifo_V_MESSAGE_29_din)           
        );
        
        initial begin
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            full = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            out_fifo_V_MESSAGE_6_din = 32'h00000008;
            out_fifo_V_MESSAGE_7_din = 32'h00000009;
            out_fifo_V_MESSAGE_8_din = 32'h0000000A;
            out_fifo_V_MESSAGE_9_din = 32'h0000000B;
            out_fifo_V_MESSAGE_10_din = 32'h0000000C;
            out_fifo_V_MESSAGE_11_din = 32'h0000000D;
            out_fifo_V_MESSAGE_12_din = 32'h0000000E;
            out_fifo_V_MESSAGE_13_din = 32'h0000000F;
            out_fifo_V_MESSAGE_14_din = 32'h00000010;
            out_fifo_V_MESSAGE_15_din = 32'h00000011;
            out_fifo_V_MESSAGE_16_din = 32'h00000012;
            out_fifo_V_MESSAGE_17_din = 32'h00000013;
            out_fifo_V_MESSAGE_18_din = 32'h00000014;
            out_fifo_V_MESSAGE_19_din = 32'h00000015;
            out_fifo_V_MESSAGE_20_din = 32'h00000016;
            out_fifo_V_MESSAGE_21_din = 32'h00000017;
            out_fifo_V_MESSAGE_22_din = 32'h00000018;
            out_fifo_V_MESSAGE_23_din = 32'h00000019;
            out_fifo_V_MESSAGE_24_din = 32'h0000001A;
            out_fifo_V_MESSAGE_25_din = 32'h0000001B;
            out_fifo_V_MESSAGE_26_din = 32'h0000001C;
            out_fifo_V_MESSAGE_27_din = 32'h0000001D;
            out_fifo_V_MESSAGE_28_din = 32'h0000001E;
            out_fifo_V_MESSAGE_29_din = 32'h0000001F;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'hFF;
            out_fifo_V_BS_ID_write = 1;
            full = 1;
            
            
            out_fifo_V_FPGA_ID_din = 8'hFF;
            out_fifo_V_PCKG_ID_din = 16'hFFFF;
            out_fifo_V_TX_UID_din = 8'hFF;
            out_fifo_V_RX_UID_din = 8'hFF;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'hFFFE;
            
            out_fifo_V_MESSAGE_0_din = 32'hFFFFFFFD;
            out_fifo_V_MESSAGE_1_din = 32'hFFFFFFFC;
            out_fifo_V_MESSAGE_2_din = 32'hFFFFFFFB;
            out_fifo_V_MESSAGE_3_din = 32'hFFFFFFFA;
            out_fifo_V_MESSAGE_4_din = 32'hFFFFFFF9;
            out_fifo_V_MESSAGE_5_din = 32'hFFFFFFF8;
            out_fifo_V_MESSAGE_6_din = 32'hFFFFFFF7;
            out_fifo_V_MESSAGE_7_din = 32'hFFFFFFF6;
            out_fifo_V_MESSAGE_8_din = 32'hFFFFFFF5;
            out_fifo_V_MESSAGE_9_din = 32'hFFFFFFF4;
            out_fifo_V_MESSAGE_10_din = 32'hFFFFFFF3;
            out_fifo_V_MESSAGE_11_din = 32'hFFFFFFF2;
            out_fifo_V_MESSAGE_12_din = 32'hFFFFFFF1;
            out_fifo_V_MESSAGE_13_din = 32'hFFFFFFF0;
            out_fifo_V_MESSAGE_14_din = 32'hFFFFFFFF;
            out_fifo_V_MESSAGE_15_din = 32'hFFFFFFEE;
            out_fifo_V_MESSAGE_16_din = 32'hFFFFFFDD;
            out_fifo_V_MESSAGE_17_din = 32'hFFFFFFCC;
            out_fifo_V_MESSAGE_18_din = 32'hFFFFFFBB;
            out_fifo_V_MESSAGE_19_din = 32'hFFFFFFAA;
            out_fifo_V_MESSAGE_20_din = 32'hFFFFFF99;
            out_fifo_V_MESSAGE_21_din = 32'hFFFFFF88;
            out_fifo_V_MESSAGE_22_din = 32'hFFFFFF77;
            out_fifo_V_MESSAGE_23_din = 32'hFFFFFF66;
            out_fifo_V_MESSAGE_24_din = 32'hFFFFFF55;
            out_fifo_V_MESSAGE_25_din = 32'hFFFFFF44;
            out_fifo_V_MESSAGE_26_din = 32'hFFFFFF33;
            out_fifo_V_MESSAGE_27_din = 32'hFFFFFF22;
            out_fifo_V_MESSAGE_28_din = 32'hFFFFFF11;
            out_fifo_V_MESSAGE_29_din = 32'hFFFFFF00;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 0;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0000;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000000;
            out_fifo_V_MESSAGE_1_din = 32'h00000000;
            out_fifo_V_MESSAGE_2_din = 32'h00000000;
            out_fifo_V_MESSAGE_3_din = 32'h00000000;
            out_fifo_V_MESSAGE_4_din = 32'h00000000;
            out_fifo_V_MESSAGE_5_din = 32'h00000000;
            out_fifo_V_MESSAGE_6_din = 32'h00000000;
            out_fifo_V_MESSAGE_7_din = 32'h00000000;
            out_fifo_V_MESSAGE_8_din = 32'h00000000;
            out_fifo_V_MESSAGE_9_din = 32'h00000000;
            out_fifo_V_MESSAGE_10_din = 32'h00000000;
            out_fifo_V_MESSAGE_11_din = 32'h00000000;
            out_fifo_V_MESSAGE_12_din = 32'h00000000;
            out_fifo_V_MESSAGE_13_din = 32'h00000000;
            out_fifo_V_MESSAGE_14_din = 32'h00000000;
            out_fifo_V_MESSAGE_15_din = 32'h00000000;
            out_fifo_V_MESSAGE_16_din = 32'h00000000;
            out_fifo_V_MESSAGE_17_din = 32'h00000000;
            out_fifo_V_MESSAGE_18_din = 32'h00000000;
            out_fifo_V_MESSAGE_19_din = 32'h00000000;
            out_fifo_V_MESSAGE_20_din = 32'h00000000;
            out_fifo_V_MESSAGE_21_din = 32'h00000000;
            out_fifo_V_MESSAGE_22_din = 32'h00000000;
            out_fifo_V_MESSAGE_23_din = 32'h00000000;
            out_fifo_V_MESSAGE_24_din = 32'h00000000;
            out_fifo_V_MESSAGE_25_din = 32'h00000000;
            out_fifo_V_MESSAGE_26_din = 32'h00000000;
            out_fifo_V_MESSAGE_27_din = 32'h00000000;
            out_fifo_V_MESSAGE_28_din = 32'h00000000;
            out_fifo_V_MESSAGE_29_din = 32'h00000000;
            
            #400;
            
            out_fifo_V_BS_ID_din = 8'h00;
            out_fifo_V_BS_ID_write = 1;
            
            out_fifo_V_FPGA_ID_din = 8'h00;
            out_fifo_V_PCKG_ID_din = 16'h0000;
            out_fifo_V_TX_UID_din = 8'h00;
            out_fifo_V_RX_UID_din = 8'h00;
            out_fifo_V_VALID_PACKET_BYTES_din = 16'h0001;
            
            out_fifo_V_MESSAGE_0_din = 32'h00000002;
            out_fifo_V_MESSAGE_1_din = 32'h00000003;
            out_fifo_V_MESSAGE_2_din = 32'h00000004;
            out_fifo_V_MESSAGE_3_din = 32'h00000005;
            out_fifo_V_MESSAGE_4_din = 32'h00000006;
            out_fifo_V_MESSAGE_5_din = 32'h00000007;
            out_fifo_V_MESSAGE_6_din = 32'h00000008;
            out_fifo_V_MESSAGE_7_din = 32'h00000009;
            out_fifo_V_MESSAGE_8_din = 32'h0000000A;
            out_fifo_V_MESSAGE_9_din = 32'h0000000B;
            out_fifo_V_MESSAGE_10_din = 32'h0000000C;
            out_fifo_V_MESSAGE_11_din = 32'h0000000D;
            out_fifo_V_MESSAGE_12_din = 32'h0000000E;
            out_fifo_V_MESSAGE_13_din = 32'h0000000F;
            out_fifo_V_MESSAGE_14_din = 32'h00000010;
            out_fifo_V_MESSAGE_15_din = 32'h00000011;
            out_fifo_V_MESSAGE_16_din = 32'h00000012;
            out_fifo_V_MESSAGE_17_din = 32'h00000013;
            out_fifo_V_MESSAGE_18_din = 32'h00000014;
            out_fifo_V_MESSAGE_19_din = 32'h00000015;
            out_fifo_V_MESSAGE_20_din = 32'h00000016;
            out_fifo_V_MESSAGE_21_din = 32'h00000017;
            out_fifo_V_MESSAGE_22_din = 32'h00000018;
            out_fifo_V_MESSAGE_23_din = 32'h00000019;
            out_fifo_V_MESSAGE_24_din = 32'h0000001A;
            out_fifo_V_MESSAGE_25_din = 32'h0000001B;
            out_fifo_V_MESSAGE_26_din = 32'h0000001C;
            out_fifo_V_MESSAGE_27_din = 32'h0000001D;
            out_fifo_V_MESSAGE_28_din = 32'h0000001E;
            out_fifo_V_MESSAGE_29_din = 32'h0000001F;
            
        end
        
    
    endmodule

`else
	// Statements
`endif 
