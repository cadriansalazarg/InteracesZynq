`timescale 1ns / 1ps

`define PACKET_SIZE_256  //Debe ajustarse al tamaño de paquete que mejor se ajusta, de manera que concuerde con PACKET_SIZE_BITS, o al menos PACKET_SIZE_BITS sea menor o igual que este parámetro
//`define PACKET_SIZE_512
//`define PACKET_SIZE_1024

`ifdef PACKET_SIZE_256
    
    module  FIFO_to_Custom_IP #(parameter PACKET_SIZE_BITS = 256)
        (
        rd_en, dout, empty, 
        in_fifo_V_BS_ID_dout, in_fifo_V_BS_ID_empty_n, in_fifo_V_BS_ID_read,
        in_fifo_V_FPGA_ID_dout, in_fifo_V_FPGA_ID_empty_n,
        in_fifo_V_PCKG_ID_dout, in_fifo_V_PCKG_ID_empty_n,
        in_fifo_V_TX_UID_dout, in_fifo_V_TX_UID_empty_n,
        in_fifo_V_RX_UID_dout, in_fifo_V_RX_UID_empty_n,
        in_fifo_V_VALID_PACKET_BYTES_dout, in_fifo_V_VALID_PACKET_BYTES_empty_n,
        in_fifo_V_MESSAGE_0_dout, in_fifo_V_MESSAGE_0_empty_n,
        in_fifo_V_MESSAGE_1_dout, in_fifo_V_MESSAGE_1_empty_n,
        in_fifo_V_MESSAGE_2_dout, in_fifo_V_MESSAGE_2_empty_n,
        in_fifo_V_MESSAGE_3_dout, in_fifo_V_MESSAGE_3_empty_n,
        in_fifo_V_MESSAGE_4_dout, in_fifo_V_MESSAGE_4_empty_n,
        in_fifo_V_MESSAGE_5_dout, in_fifo_V_MESSAGE_5_empty_n
        );
        
        
        input [PACKET_SIZE_BITS-1:0] dout;
        input empty;
        output rd_en;
        
        output [7:0] in_fifo_V_BS_ID_dout;
        output in_fifo_V_BS_ID_empty_n;
        input in_fifo_V_BS_ID_read;
        
        output [7:0] in_fifo_V_FPGA_ID_dout;
        output in_fifo_V_FPGA_ID_empty_n;
        
        output [15:0] in_fifo_V_PCKG_ID_dout;
        output in_fifo_V_PCKG_ID_empty_n;
        
        output [7:0] in_fifo_V_TX_UID_dout;
        output in_fifo_V_TX_UID_empty_n;
        
        output [7:0] in_fifo_V_RX_UID_dout;
        output in_fifo_V_RX_UID_empty_n;
        
        output [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        output in_fifo_V_VALID_PACKET_BYTES_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_0_dout;
        output in_fifo_V_MESSAGE_0_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_1_dout;
        output in_fifo_V_MESSAGE_1_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_2_dout;
        output in_fifo_V_MESSAGE_2_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_3_dout;
        output in_fifo_V_MESSAGE_3_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_4_dout;
        output in_fifo_V_MESSAGE_4_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_5_dout;
        output in_fifo_V_MESSAGE_5_empty_n;
        
        wire not_empty;
        assign not_empty = ~empty;
        
        
        assign rd_en = in_fifo_V_BS_ID_read;
        assign in_fifo_V_BS_ID_dout = dout[255:248];
        assign in_fifo_V_BS_ID_empty_n = not_empty;
        assign in_fifo_V_FPGA_ID_dout = dout[247:240];
        assign in_fifo_V_FPGA_ID_empty_n = not_empty;
        assign in_fifo_V_PCKG_ID_dout = dout[239:224];
        assign in_fifo_V_PCKG_ID_empty_n = not_empty;
        assign in_fifo_V_TX_UID_dout = dout[223:216];
        assign in_fifo_V_TX_UID_empty_n = not_empty;
        assign in_fifo_V_RX_UID_dout = dout[215:208];
        assign in_fifo_V_RX_UID_empty_n = not_empty;
        assign in_fifo_V_VALID_PACKET_BYTES_dout = dout[207:192];
        assign in_fifo_V_VALID_PACKET_BYTES_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_0_dout = dout[191:160];
        assign in_fifo_V_MESSAGE_0_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_1_dout = dout[159:128];
        assign in_fifo_V_MESSAGE_1_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_2_dout = dout[127:96];
        assign in_fifo_V_MESSAGE_2_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_3_dout = dout[95:64];
        assign in_fifo_V_MESSAGE_3_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_4_dout = dout[63:32];
        assign in_fifo_V_MESSAGE_4_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_5_dout = dout[31:0];
        assign in_fifo_V_MESSAGE_5_empty_n = not_empty;
         
    endmodule 
           
`elsif PACKET_SIZE_512

    module  FIFO_to_Custom_IP #(parameter PACKET_SIZE_BITS = 512)
        (
        rd_en, dout, empty, 
        in_fifo_V_BS_ID_dout, in_fifo_V_BS_ID_empty_n, in_fifo_V_BS_ID_read,
        in_fifo_V_FPGA_ID_dout, in_fifo_V_FPGA_ID_empty_n,
        in_fifo_V_PCKG_ID_dout, in_fifo_V_PCKG_ID_empty_n,
        in_fifo_V_TX_UID_dout, in_fifo_V_TX_UID_empty_n,
        in_fifo_V_RX_UID_dout, in_fifo_V_RX_UID_empty_n,
        in_fifo_V_VALID_PACKET_BYTES_dout, in_fifo_V_VALID_PACKET_BYTES_empty_n,
        in_fifo_V_MESSAGE_0_dout, in_fifo_V_MESSAGE_0_empty_n,
        in_fifo_V_MESSAGE_1_dout, in_fifo_V_MESSAGE_1_empty_n,
        in_fifo_V_MESSAGE_2_dout, in_fifo_V_MESSAGE_2_empty_n,
        in_fifo_V_MESSAGE_3_dout, in_fifo_V_MESSAGE_3_empty_n,
        in_fifo_V_MESSAGE_4_dout, in_fifo_V_MESSAGE_4_empty_n,
        in_fifo_V_MESSAGE_5_dout, in_fifo_V_MESSAGE_5_empty_n,
        in_fifo_V_MESSAGE_6_dout, in_fifo_V_MESSAGE_6_empty_n,
        in_fifo_V_MESSAGE_7_dout, in_fifo_V_MESSAGE_7_empty_n,
        in_fifo_V_MESSAGE_8_dout, in_fifo_V_MESSAGE_8_empty_n,
        in_fifo_V_MESSAGE_9_dout, in_fifo_V_MESSAGE_9_empty_n,
        in_fifo_V_MESSAGE_10_dout, in_fifo_V_MESSAGE_10_empty_n,
        in_fifo_V_MESSAGE_11_dout, in_fifo_V_MESSAGE_11_empty_n,
        in_fifo_V_MESSAGE_12_dout, in_fifo_V_MESSAGE_12_empty_n,
        in_fifo_V_MESSAGE_13_dout, in_fifo_V_MESSAGE_13_empty_n
        );
        
        input [PACKET_SIZE_BITS-1:0] dout;
        input empty;
        output rd_en;
        
        output [7:0] in_fifo_V_BS_ID_dout;
        output in_fifo_V_BS_ID_empty_n;
        input in_fifo_V_BS_ID_read;
        
        output [7:0] in_fifo_V_FPGA_ID_dout;
        output in_fifo_V_FPGA_ID_empty_n;
        
        output [15:0] in_fifo_V_PCKG_ID_dout;
        output in_fifo_V_PCKG_ID_empty_n;
        
        output [7:0] in_fifo_V_TX_UID_dout;
        output in_fifo_V_TX_UID_empty_n;
        
        output [7:0] in_fifo_V_RX_UID_dout;
        output in_fifo_V_RX_UID_empty_n;
        
        output [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        output in_fifo_V_VALID_PACKET_BYTES_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_0_dout;
        output in_fifo_V_MESSAGE_0_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_1_dout;
        output in_fifo_V_MESSAGE_1_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_2_dout;
        output in_fifo_V_MESSAGE_2_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_3_dout;
        output in_fifo_V_MESSAGE_3_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_4_dout;
        output in_fifo_V_MESSAGE_4_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_5_dout;
        output in_fifo_V_MESSAGE_5_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_6_dout;
        output in_fifo_V_MESSAGE_6_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_7_dout;
        output in_fifo_V_MESSAGE_7_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_8_dout;
        output in_fifo_V_MESSAGE_8_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_9_dout;
        output in_fifo_V_MESSAGE_9_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_10_dout;
        output in_fifo_V_MESSAGE_10_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_11_dout;
        output in_fifo_V_MESSAGE_11_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_12_dout;
        output in_fifo_V_MESSAGE_12_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_13_dout;
        output in_fifo_V_MESSAGE_13_empty_n;
        
        wire not_empty;
        assign not_empty = ~empty;
        
        assign rd_en = in_fifo_V_BS_ID_read;
        assign in_fifo_V_BS_ID_dout = dout[511:504];
        assign in_fifo_V_BS_ID_empty_n = not_empty;
        assign in_fifo_V_FPGA_ID_dout = dout[503:496];
        assign in_fifo_V_FPGA_ID_empty_n = not_empty;
        assign in_fifo_V_PCKG_ID_dout = dout[495:480];
        assign in_fifo_V_PCKG_ID_empty_n = not_empty;
        assign in_fifo_V_TX_UID_dout = dout[479:472];
        assign in_fifo_V_TX_UID_empty_n = not_empty;
        assign in_fifo_V_RX_UID_dout = dout[471:464];
        assign in_fifo_V_RX_UID_empty_n = not_empty;
        assign in_fifo_V_VALID_PACKET_BYTES_dout = dout[463:448];
        assign in_fifo_V_VALID_PACKET_BYTES_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_0_dout = dout[447:416];
        assign in_fifo_V_MESSAGE_0_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_1_dout = dout[415:384];
        assign in_fifo_V_MESSAGE_1_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_2_dout = dout[383:352];
        assign in_fifo_V_MESSAGE_2_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_3_dout = dout[351:320];
        assign in_fifo_V_MESSAGE_3_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_4_dout = dout[319:288];
        assign in_fifo_V_MESSAGE_4_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_5_dout = dout[287:256];
        assign in_fifo_V_MESSAGE_5_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_6_dout = dout[255:224];
        assign in_fifo_V_MESSAGE_6_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_7_dout = dout[223:192];
        assign in_fifo_V_MESSAGE_7_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_8_dout = dout[191:160];
        assign in_fifo_V_MESSAGE_8_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_9_dout = dout[159:128];
        assign in_fifo_V_MESSAGE_9_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_10_dout = dout[127:96];
        assign in_fifo_V_MESSAGE_10_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_11_dout = dout[95:64];
        assign in_fifo_V_MESSAGE_11_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_12_dout = dout[63:32];
        assign in_fifo_V_MESSAGE_12_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_13_dout = dout[31:0];
        assign in_fifo_V_MESSAGE_13_empty_n = not_empty;
        
    endmodule        
 
`elsif PACKET_SIZE_1024  

    module  FIFO_to_Custom_IP #(parameter PACKET_SIZE_BITS = 1024)
        (
        rd_en, dout, empty, 
        in_fifo_V_BS_ID_dout, in_fifo_V_BS_ID_empty_n, in_fifo_V_BS_ID_read,
        in_fifo_V_FPGA_ID_dout, in_fifo_V_FPGA_ID_empty_n,
        in_fifo_V_PCKG_ID_dout, in_fifo_V_PCKG_ID_empty_n,
        in_fifo_V_TX_UID_dout, in_fifo_V_TX_UID_empty_n,
        in_fifo_V_RX_UID_dout, in_fifo_V_RX_UID_empty_n,
        in_fifo_V_VALID_PACKET_BYTES_dout, in_fifo_V_VALID_PACKET_BYTES_empty_n,
        in_fifo_V_MESSAGE_0_dout, in_fifo_V_MESSAGE_0_empty_n,
        in_fifo_V_MESSAGE_1_dout, in_fifo_V_MESSAGE_1_empty_n,
        in_fifo_V_MESSAGE_2_dout, in_fifo_V_MESSAGE_2_empty_n,
        in_fifo_V_MESSAGE_3_dout, in_fifo_V_MESSAGE_3_empty_n,
        in_fifo_V_MESSAGE_4_dout, in_fifo_V_MESSAGE_4_empty_n,
        in_fifo_V_MESSAGE_5_dout, in_fifo_V_MESSAGE_5_empty_n,
        in_fifo_V_MESSAGE_6_dout, in_fifo_V_MESSAGE_6_empty_n,
        in_fifo_V_MESSAGE_7_dout, in_fifo_V_MESSAGE_7_empty_n,
        in_fifo_V_MESSAGE_8_dout, in_fifo_V_MESSAGE_8_empty_n,
        in_fifo_V_MESSAGE_9_dout, in_fifo_V_MESSAGE_9_empty_n,
        in_fifo_V_MESSAGE_10_dout, in_fifo_V_MESSAGE_10_empty_n,
        in_fifo_V_MESSAGE_11_dout, in_fifo_V_MESSAGE_11_empty_n,
        in_fifo_V_MESSAGE_12_dout, in_fifo_V_MESSAGE_12_empty_n,
        in_fifo_V_MESSAGE_13_dout, in_fifo_V_MESSAGE_13_empty_n,
        in_fifo_V_MESSAGE_14_dout, in_fifo_V_MESSAGE_14_empty_n,
        in_fifo_V_MESSAGE_15_dout, in_fifo_V_MESSAGE_15_empty_n,
        in_fifo_V_MESSAGE_16_dout, in_fifo_V_MESSAGE_16_empty_n,
        in_fifo_V_MESSAGE_17_dout, in_fifo_V_MESSAGE_17_empty_n,
        in_fifo_V_MESSAGE_18_dout, in_fifo_V_MESSAGE_18_empty_n,
        in_fifo_V_MESSAGE_19_dout, in_fifo_V_MESSAGE_19_empty_n,
        in_fifo_V_MESSAGE_20_dout, in_fifo_V_MESSAGE_20_empty_n,
        in_fifo_V_MESSAGE_21_dout, in_fifo_V_MESSAGE_21_empty_n,
        in_fifo_V_MESSAGE_22_dout, in_fifo_V_MESSAGE_22_empty_n,
        in_fifo_V_MESSAGE_23_dout, in_fifo_V_MESSAGE_23_empty_n,
        in_fifo_V_MESSAGE_24_dout, in_fifo_V_MESSAGE_24_empty_n,
        in_fifo_V_MESSAGE_25_dout, in_fifo_V_MESSAGE_25_empty_n,
        in_fifo_V_MESSAGE_26_dout, in_fifo_V_MESSAGE_26_empty_n,
        in_fifo_V_MESSAGE_27_dout, in_fifo_V_MESSAGE_27_empty_n,
        in_fifo_V_MESSAGE_28_dout, in_fifo_V_MESSAGE_28_empty_n,
        in_fifo_V_MESSAGE_29_dout, in_fifo_V_MESSAGE_29_empty_n
        );
        
        input [PACKET_SIZE_BITS-1:0] dout;
        input empty;
        output rd_en;
        
        output [7:0] in_fifo_V_BS_ID_dout;
        output in_fifo_V_BS_ID_empty_n;
        input in_fifo_V_BS_ID_read;
        
        output [7:0] in_fifo_V_FPGA_ID_dout;
        output in_fifo_V_FPGA_ID_empty_n;
        
        output [15:0] in_fifo_V_PCKG_ID_dout;
        output in_fifo_V_PCKG_ID_empty_n;
        
        output [7:0] in_fifo_V_TX_UID_dout;
        output in_fifo_V_TX_UID_empty_n;
        
        output [7:0] in_fifo_V_RX_UID_dout;
        output in_fifo_V_RX_UID_empty_n;
        
        output [15:0] in_fifo_V_VALID_PACKET_BYTES_dout;
        output in_fifo_V_VALID_PACKET_BYTES_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_0_dout;
        output in_fifo_V_MESSAGE_0_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_1_dout;
        output in_fifo_V_MESSAGE_1_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_2_dout;
        output in_fifo_V_MESSAGE_2_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_3_dout;
        output in_fifo_V_MESSAGE_3_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_4_dout;
        output in_fifo_V_MESSAGE_4_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_5_dout;
        output in_fifo_V_MESSAGE_5_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_6_dout;
        output in_fifo_V_MESSAGE_6_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_7_dout;
        output in_fifo_V_MESSAGE_7_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_8_dout;
        output in_fifo_V_MESSAGE_8_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_9_dout;
        output in_fifo_V_MESSAGE_9_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_10_dout;
        output in_fifo_V_MESSAGE_10_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_11_dout;
        output in_fifo_V_MESSAGE_11_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_12_dout;
        output in_fifo_V_MESSAGE_12_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_13_dout;
        output in_fifo_V_MESSAGE_13_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_14_dout;
        output in_fifo_V_MESSAGE_14_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_15_dout;
        output in_fifo_V_MESSAGE_15_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_16_dout;
        output in_fifo_V_MESSAGE_16_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_17_dout;
        output in_fifo_V_MESSAGE_17_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_18_dout;
        output in_fifo_V_MESSAGE_18_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_19_dout;
        output in_fifo_V_MESSAGE_19_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_20_dout;
        output in_fifo_V_MESSAGE_20_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_21_dout;
        output in_fifo_V_MESSAGE_21_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_22_dout;
        output in_fifo_V_MESSAGE_22_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_23_dout;
        output in_fifo_V_MESSAGE_23_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_24_dout;
        output in_fifo_V_MESSAGE_24_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_25_dout;
        output in_fifo_V_MESSAGE_25_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_26_dout;
        output in_fifo_V_MESSAGE_26_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_27_dout;
        output in_fifo_V_MESSAGE_27_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_28_dout;
        output in_fifo_V_MESSAGE_28_empty_n;
        
        output [31:0] in_fifo_V_MESSAGE_29_dout;
        output in_fifo_V_MESSAGE_29_empty_n;
        
        wire not_empty;
        assign not_empty = ~empty;
        
        assign rd_en = in_fifo_V_BS_ID_read;
        assign in_fifo_V_BS_ID_dout = dout[1023:1016];
        assign in_fifo_V_BS_ID_empty_n = not_empty;
        assign in_fifo_V_FPGA_ID_dout = dout[1015:1008];
        assign in_fifo_V_FPGA_ID_empty_n = not_empty;
        assign in_fifo_V_PCKG_ID_dout = dout[1007:992];
        assign in_fifo_V_PCKG_ID_empty_n = not_empty;
        assign in_fifo_V_TX_UID_dout = dout[991:984];
        assign in_fifo_V_TX_UID_empty_n = not_empty;
        assign in_fifo_V_RX_UID_dout = dout[983:976];
        assign in_fifo_V_RX_UID_empty_n = not_empty;
        assign in_fifo_V_VALID_PACKET_BYTES_dout = dout[975:960];
        assign in_fifo_V_VALID_PACKET_BYTES_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_0_dout = dout[959:928];
        assign in_fifo_V_MESSAGE_0_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_1_dout = dout[927:896];
        assign in_fifo_V_MESSAGE_1_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_2_dout = dout[895:864];
        assign in_fifo_V_MESSAGE_2_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_3_dout = dout[863:832];
        assign in_fifo_V_MESSAGE_3_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_4_dout = dout[831:800];
        assign in_fifo_V_MESSAGE_4_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_5_dout = dout[799:768];
        assign in_fifo_V_MESSAGE_5_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_6_dout = dout[767:736];
        assign in_fifo_V_MESSAGE_6_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_7_dout = dout[735:704];
        assign in_fifo_V_MESSAGE_7_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_8_dout = dout[703:672];
        assign in_fifo_V_MESSAGE_8_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_9_dout = dout[671:640];
        assign in_fifo_V_MESSAGE_9_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_10_dout = dout[639:608];
        assign in_fifo_V_MESSAGE_10_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_11_dout = dout[607:576];
        assign in_fifo_V_MESSAGE_11_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_12_dout = dout[575:544];
        assign in_fifo_V_MESSAGE_12_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_13_dout = dout[543:512];
        assign in_fifo_V_MESSAGE_13_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_14_dout = dout[511:490];
        assign in_fifo_V_MESSAGE_14_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_15_dout = dout[479:448];
        assign in_fifo_V_MESSAGE_15_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_16_dout = dout[447:416];
        assign in_fifo_V_MESSAGE_16_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_17_dout = dout[415:384];
        assign in_fifo_V_MESSAGE_17_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_18_dout = dout[383:352];
        assign in_fifo_V_MESSAGE_18_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_19_dout = dout[351:320];
        assign in_fifo_V_MESSAGE_19_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_20_dout = dout[319:288];
        assign in_fifo_V_MESSAGE_20_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_21_dout = dout[287:256];
        assign in_fifo_V_MESSAGE_21_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_22_dout = dout[255:224];
        assign in_fifo_V_MESSAGE_22_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_23_dout = dout[223:192];
        assign in_fifo_V_MESSAGE_23_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_24_dout = dout[191:160];
        assign in_fifo_V_MESSAGE_24_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_25_dout = dout[159:128];
        assign in_fifo_V_MESSAGE_25_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_26_dout = dout[127:96];
        assign in_fifo_V_MESSAGE_26_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_27_dout = dout[95:64];
        assign in_fifo_V_MESSAGE_27_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_28_dout = dout[63:32];
        assign in_fifo_V_MESSAGE_28_empty_n = not_empty;
        assign in_fifo_V_MESSAGE_29_dout = dout[31:0];
        assign in_fifo_V_MESSAGE_29_empty_n = not_empty;
        
        
    endmodule     
 
`else
	// Statements
`endif   
    

