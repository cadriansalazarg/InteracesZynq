`timescale 1ns / 1ps

`define PACKET_SIZE_128

module register #(parameter WIDTH = 32) (user_clk, RST, Enable, D, Q);

	output reg [WIDTH-1: 0] Q;
	input user_clk, RST, Enable;
	input [WIDTH-1: 0] D;
	
	always @(posedge user_clk)
      if (RST) begin
         Q <= 0;
      end else if (Enable) begin
         Q <= D;
      end
endmodule 

module ROM (CLK, Address, Output);
	
	input CLK;
	input [7:0] Address;  // TX_UID
	output reg [7:0] Output;  // BUS_ID
   
   always @(posedge CLK)
		case (Address)
			8'b00000000: Output <= 8'b00000000;
         8'b00000001: Output <= 8'b00000011;
         8'b00000010: Output <= 8'b00000000;
         8'b00000011: Output <= 8'b00000000;
         8'b00000100: Output <= 8'b00000000;
         8'b00000101: Output <= 8'b00000000;
         8'b00000110: Output <= 8'b00000000;
         8'b00000111: Output <= 8'b00000000;
         8'b00001000: Output <= 8'b00000000;
         8'b00001001: Output <= 8'b00000000;
         8'b00001010: Output <= 8'b00000000;
         8'b00001011: Output <= 8'b00000000;
         8'b00001100: Output <= 8'b00000000;
         8'b00001101: Output <= 8'b00000000;
         8'b00001110: Output <= 8'b00000000;
         8'b00001111: Output <= 8'b00000000;
         default: Output <= 8'b11111111;
     endcase
endmodule


module receiver #(parameter PACKET_SIZE = 128, RX_TDATA_SIZE = 32) 
(user_clk, RST, start, din, wr_en, full, m_axi_rx_tdata, m_axi_rx_tlast, m_axi_rx_tvalid, Error);
	
	localparam NUMBER_OF_PACKETS = PACKET_SIZE/RX_TDATA_SIZE;
	
	localparam S0 = 3'd0, S1 = 3'd1, S2 = 3'd2, S3 = 3'd3, S4 = 3'd4, S5 = 3'd5, S6 = 3'd6, S7 = 3'd7;
	reg [2:0] State, NextState;
	
	input user_clk, RST, start;
	
	output [PACKET_SIZE-1:0]  din ;
	output reg wr_en;
	input full;
	output reg Error;
	
	input [RX_TDATA_SIZE-1:0] m_axi_rx_tdata;
	input m_axi_rx_tlast, m_axi_rx_tvalid;
	
	wire [PACKET_SIZE-1:0]  din_reg ;
	wire [7:0] BS_ID;
	
	reg  m_axi_rx_tlast_reg, m_axi_rx_tvalid_reg;
	reg start_reg;
	reg [RX_TDATA_SIZE-1:0] m_axi_rx_tdata_reg;
	reg [RX_TDATA_SIZE-1:0] m_axi_rx_tdata_reg1;
	reg full_reg;
	reg reset_output_register, wr_en_reg, reset_file_register, enable_output_register;
	
	reg [7:0] Q_seq_counter;
	
	// **************** Parallel Register ********************************************************************
	
	always @(posedge user_clk)
		if (RST) begin 
			m_axi_rx_tlast_reg <= 1'b0;
			m_axi_rx_tvalid_reg <= 1'b0;
			m_axi_rx_tdata_reg <= 0;
			start_reg <= 0;
			full_reg <= 0;
			wr_en <= 0;
		end else begin
			m_axi_rx_tlast_reg <= m_axi_rx_tlast;
			m_axi_rx_tvalid_reg <= m_axi_rx_tvalid;
			m_axi_rx_tdata_reg <= m_axi_rx_tdata;
			start_reg <= start;
			full_reg <= full;
			wr_en <= wr_en_reg;
		end
		
	always @(posedge user_clk)
		if (RST  | reset_file_register) begin 
			m_axi_rx_tdata_reg1 <= 0;
		end else if (m_axi_rx_tvalid_reg) begin
			m_axi_rx_tdata_reg1 <= m_axi_rx_tdata_reg;
		end


// *********************************** Counter and decoder in function of packet size ********************************
`ifdef PACKET_SIZE_4096
	reg [6:0] Q_counter;
	reg [127:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				7'd0  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
				7'd1  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
				7'd2  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
				7'd3  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
				7'd4  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
				7'd5  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
				7'd6  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
				7'd7  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
				7'd8  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
				7'd9  : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
				7'd10 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
				7'd11 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
				7'd12 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
				7'd13 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
				7'd14 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
				7'd15 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;	
				7'd16 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
				7'd17 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
				7'd18 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
				7'd19 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
				7'd20 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
				7'd21 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
				7'd22 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
				7'd23 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
				7'd24 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
				7'd25 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
				7'd26 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
				7'd27 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
				7'd28 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
				7'd29 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
				7'd30 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
				7'd31 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
				7'd32 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
				7'd33 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
				7'd34 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
				7'd35 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
				7'd36 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
				7'd37 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
				7'd38 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
				7'd39 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
				7'd40 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
				7'd41 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
				7'd42 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
				7'd43 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
				7'd44 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
				7'd45 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
				7'd46 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
				7'd47 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;	
				7'd48 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
				7'd49 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
				7'd50 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
				7'd51 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
				7'd52 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
				7'd53 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
				7'd54 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
				7'd55 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
				7'd56 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
				7'd57 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
				7'd58 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
				7'd59 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
				7'd60 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
				7'd61 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
				7'd62 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
				7'd63 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
				7'd64 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
				7'd65 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
				7'd66 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
				7'd67 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
				7'd68 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
				7'd69 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
				7'd70 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
				7'd71 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
				7'd72 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd73 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd74 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd75 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd76 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd77 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd78 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd79 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;	
				7'd80 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd81 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd82 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd83 : Enable_Registers <= 128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd84 : Enable_Registers <= 128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd85 : Enable_Registers <= 128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd86 : Enable_Registers <= 128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd87 : Enable_Registers <= 128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd88 : Enable_Registers <= 128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd89 : Enable_Registers <= 128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd90 : Enable_Registers <= 128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd91 : Enable_Registers <= 128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd92 : Enable_Registers <= 128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd93 : Enable_Registers <= 128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd94 : Enable_Registers <= 128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd95 : Enable_Registers <= 128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd96 : Enable_Registers <= 128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd97 : Enable_Registers <= 128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd98 : Enable_Registers <= 128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd99 : Enable_Registers <= 128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd100: Enable_Registers <= 128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd101: Enable_Registers <= 128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd102: Enable_Registers <= 128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd103: Enable_Registers <= 128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd104: Enable_Registers <= 128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd105: Enable_Registers <= 128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd106: Enable_Registers <= 128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd107: Enable_Registers <= 128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd108: Enable_Registers <= 128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd109: Enable_Registers <= 128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd110: Enable_Registers <= 128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd111: Enable_Registers <= 128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;	
				7'd112: Enable_Registers <= 128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd113: Enable_Registers <= 128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd114: Enable_Registers <= 128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd115: Enable_Registers <= 128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd116: Enable_Registers <= 128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd117: Enable_Registers <= 128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd118: Enable_Registers <= 128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd119: Enable_Registers <= 128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd120: Enable_Registers <= 128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd121: Enable_Registers <= 128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd122: Enable_Registers <= 128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd123: Enable_Registers <= 128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd124: Enable_Registers <= 128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd125: Enable_Registers <= 128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd126: Enable_Registers <= 128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				7'd127: Enable_Registers <= 128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_2048
	reg [5:0] Q_counter;
	reg [63:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				6'd0  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
				6'd1  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
				6'd2  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
				6'd3  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
				6'd4  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
				6'd5  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
				6'd6  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
				6'd7  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
				6'd8  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
				6'd9  : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000001000000000;
				6'd10 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000010000000000;
				6'd11 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000000100000000000;
				6'd12 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000001000000000000;
				6'd13 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000010000000000000;
				6'd14 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000000100000000000000;
				6'd15 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000001000000000000000;	
				6'd16 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000010000000000000000;
				6'd17 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000000100000000000000000;
				6'd18 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
				6'd19 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000010000000000000000000;
				6'd20 : Enable_Registers <= 64'b0000000000000000000000000000000000000000000100000000000000000000;
				6'd21 : Enable_Registers <= 64'b0000000000000000000000000000000000000000001000000000000000000000;
				6'd22 : Enable_Registers <= 64'b0000000000000000000000000000000000000000010000000000000000000000;
				6'd23 : Enable_Registers <= 64'b0000000000000000000000000000000000000000100000000000000000000000;
				6'd24 : Enable_Registers <= 64'b0000000000000000000000000000000000000001000000000000000000000000;
				6'd25 : Enable_Registers <= 64'b0000000000000000000000000000000000000010000000000000000000000000;
				6'd26 : Enable_Registers <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
				6'd27 : Enable_Registers <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
				6'd28 : Enable_Registers <= 64'b0000000000000000000000000000000000010000000000000000000000000000;
				6'd29 : Enable_Registers <= 64'b0000000000000000000000000000000000100000000000000000000000000000;
				6'd30 : Enable_Registers <= 64'b0000000000000000000000000000000001000000000000000000000000000000;
				6'd31 : Enable_Registers <= 64'b0000000000000000000000000000000010000000000000000000000000000000;
				6'd32 : Enable_Registers <= 64'b0000000000000000000000000000000100000000000000000000000000000000;
				6'd33 : Enable_Registers <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
				6'd34 : Enable_Registers <= 64'b0000000000000000000000000000010000000000000000000000000000000000;
				6'd35 : Enable_Registers <= 64'b0000000000000000000000000000100000000000000000000000000000000000;
				6'd36 : Enable_Registers <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
				6'd37 : Enable_Registers <= 64'b0000000000000000000000000010000000000000000000000000000000000000;
				6'd38 : Enable_Registers <= 64'b0000000000000000000000000100000000000000000000000000000000000000;
				6'd39 : Enable_Registers <= 64'b0000000000000000000000001000000000000000000000000000000000000000;
				6'd40 : Enable_Registers <= 64'b0000000000000000000000010000000000000000000000000000000000000000;
				6'd41 : Enable_Registers <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
				6'd42 : Enable_Registers <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
				6'd43 : Enable_Registers <= 64'b0000000000000000000010000000000000000000000000000000000000000000;
				6'd44 : Enable_Registers <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
				6'd45 : Enable_Registers <= 64'b0000000000000000001000000000000000000000000000000000000000000000;
				6'd46 : Enable_Registers <= 64'b0000000000000000010000000000000000000000000000000000000000000000;
				6'd47 : Enable_Registers <= 64'b0000000000000000100000000000000000000000000000000000000000000000;	
				6'd48 : Enable_Registers <= 64'b0000000000000001000000000000000000000000000000000000000000000000;
				6'd49 : Enable_Registers <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
				6'd50 : Enable_Registers <= 64'b0000000000000100000000000000000000000000000000000000000000000000;
				6'd51 : Enable_Registers <= 64'b0000000000001000000000000000000000000000000000000000000000000000;
				6'd52 : Enable_Registers <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
				6'd53 : Enable_Registers <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
				6'd54 : Enable_Registers <= 64'b0000000001000000000000000000000000000000000000000000000000000000;
				6'd55 : Enable_Registers <= 64'b0000000010000000000000000000000000000000000000000000000000000000;
				6'd56 : Enable_Registers <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
				6'd57 : Enable_Registers <= 64'b0000001000000000000000000000000000000000000000000000000000000000;
				6'd58 : Enable_Registers <= 64'b0000010000000000000000000000000000000000000000000000000000000000;
				6'd59 : Enable_Registers <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
				6'd60 : Enable_Registers <= 64'b0001000000000000000000000000000000000000000000000000000000000000;
				6'd61 : Enable_Registers <= 64'b0010000000000000000000000000000000000000000000000000000000000000;
				6'd62 : Enable_Registers <= 64'b0100000000000000000000000000000000000000000000000000000000000000;
				6'd63 : Enable_Registers <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_1024
	reg [4:0] Q_counter;
	reg [31:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				5'd0  : Enable_Registers <= 32'b00000000000000000000000000000001;
				5'd1  : Enable_Registers <= 32'b00000000000000000000000000000010;
				5'd2  : Enable_Registers <= 32'b00000000000000000000000000000100;
				5'd3  : Enable_Registers <= 32'b00000000000000000000000000001000;
				5'd4  : Enable_Registers <= 32'b00000000000000000000000000010000;
				5'd5  : Enable_Registers <= 32'b00000000000000000000000000100000;
				5'd6  : Enable_Registers <= 32'b00000000000000000000000001000000;
				5'd7  : Enable_Registers <= 32'b00000000000000000000000010000000;
				5'd8  : Enable_Registers <= 32'b00000000000000000000000100000000;
				5'd9  : Enable_Registers <= 32'b00000000000000000000001000000000;
				5'd10 : Enable_Registers <= 32'b00000000000000000000010000000000;
				5'd11 : Enable_Registers <= 32'b00000000000000000000100000000000;
				5'd12 : Enable_Registers <= 32'b00000000000000000001000000000000;
				5'd13 : Enable_Registers <= 32'b00000000000000000010000000000000;
				5'd14 : Enable_Registers <= 32'b00000000000000000100000000000000;
				5'd15 : Enable_Registers <= 32'b00000000000000001000000000000000;	
				5'd16 : Enable_Registers <= 32'b00000000000000010000000000000000;
				5'd17 : Enable_Registers <= 32'b00000000000000100000000000000000;
				5'd18 : Enable_Registers <= 32'b00000000000001000000000000000000;
				5'd19 : Enable_Registers <= 32'b00000000000010000000000000000000;
				5'd20 : Enable_Registers <= 32'b00000000000100000000000000000000;
				5'd21 : Enable_Registers <= 32'b00000000001000000000000000000000;
				5'd22 : Enable_Registers <= 32'b00000000010000000000000000000000;
				5'd23 : Enable_Registers <= 32'b00000000100000000000000000000000;
				5'd24 : Enable_Registers <= 32'b00000001000000000000000000000000;
				5'd25 : Enable_Registers <= 32'b00000010000000000000000000000000;
				5'd26 : Enable_Registers <= 32'b00000100000000000000000000000000;
				5'd27 : Enable_Registers <= 32'b00001000000000000000000000000000;
				5'd28 : Enable_Registers <= 32'b00010000000000000000000000000000;
				5'd29 : Enable_Registers <= 32'b00100000000000000000000000000000;
				5'd30 : Enable_Registers <= 32'b01000000000000000000000000000000;
				5'd31 : Enable_Registers <= 32'b10000000000000000000000000000000;
			endcase
`elsif PACKET_SIZE_512
	reg [3:0] Q_counter;
	reg [15:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				4'd0  : Enable_Registers <= 16'b0000000000000001;
				4'd1  : Enable_Registers <= 16'b0000000000000010;
				4'd2  : Enable_Registers <= 16'b0000000000000100;
				4'd3  : Enable_Registers <= 16'b0000000000001000;
				4'd4  : Enable_Registers <= 16'b0000000000010000;
				4'd5  : Enable_Registers <= 16'b0000000000100000;
				4'd6  : Enable_Registers <= 16'b0000000001000000;
				4'd7  : Enable_Registers <= 16'b0000000010000000;
				4'd8  : Enable_Registers <= 16'b0000000100000000;
				4'd9  : Enable_Registers <= 16'b0000001000000000;
				4'd10 : Enable_Registers <= 16'b0000010000000000;
				4'd11 : Enable_Registers <= 16'b0000100000000000;
				4'd12 : Enable_Registers <= 16'b0001000000000000;
				4'd13 : Enable_Registers <= 16'b0010000000000000;
				4'd14 : Enable_Registers <= 16'b0100000000000000;
				4'd15 : Enable_Registers <= 16'b1000000000000000;	
			endcase
`elsif PACKET_SIZE_256
	reg [2:0] Q_counter;
	reg [7:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter | reset_file_register)
				3'd0  : Enable_Registers <= 8'b00000001;
				3'd1  : Enable_Registers <= 8'b00000010;
				3'd2  : Enable_Registers <= 8'b00000100;
				3'd3  : Enable_Registers <= 8'b00001000;
				3'd4  : Enable_Registers <= 8'b00010000;
				3'd5  : Enable_Registers <= 8'b00100000;
				3'd6  : Enable_Registers <= 8'b01000000;
				3'd7  : Enable_Registers <= 8'b10000000;
			endcase
`elsif PACKET_SIZE_128
	reg [1:0] Q_counter;
	reg [3:0] Enable_Registers;
		
   always @(posedge user_clk)
      if (RST | reset_file_register)
         Q_counter <= 0;
      else if (m_axi_rx_tvalid_reg)
            Q_counter <= Q_counter + 1'b1;
				
	always @(posedge user_clk)
		if (RST | reset_file_register)	
			 Enable_Registers <= 0;
		else 
			case (Q_counter)
				2'd0  : Enable_Registers <= 4'b0001;
				2'd1  : Enable_Registers <= 4'b0010;
				2'd2  : Enable_Registers <= 4'b0100;
				2'd3  : Enable_Registers <= 4'b1000;
			endcase
`else
	// Statements
`endif


	
	
	
	// Declare a temporary loop variable to be used during
	// generation and won't be available during simulation
	genvar i;

	// Generate for loop to instantiate N times
	generate
		for (i = 0; i < NUMBER_OF_PACKETS; i = i + 1) begin : Register_Bank
          register #(.WIDTH(RX_TDATA_SIZE)) u0 (.user_clk(user_clk), .RST(RST), .Enable(Enable_Registers[i]), .D(m_axi_rx_tdata_reg1), .Q(din_reg[ (((32*NUMBER_OF_PACKETS)-1)-(i*32)) :  (((32*NUMBER_OF_PACKETS)-32)-(i*32)) ]));
		end
	endgenerate
	
	
	// ******************************************************  FSM *************************************************
	
	// Registro de estado
	always @(posedge user_clk) begin
	    if(RST)
	        State<=S0;
	    else
	        State<=NextState;
	end
	
	// L�gica combinacional de estado siguiente
	always @* begin
	    case(State)
	        S0: begin  // Wait for start providing for initialization module
                if (start_reg) NextState <= S1;
            	 else NextState <= S0;
				end
				S1: begin // Wait for tlast               // Reset output register
                if (m_axi_rx_tlast_reg) NextState <= S2;
            	 else NextState <= S1;
				end
				S2: begin // Wait for one clock cycle, for writing the last register in the register bank
                NextState <= S3;
				end
				S3: begin // Load output register and reset all the register file and counter
					 NextState <= S4;
            end	
				S4: begin // Wait if fifo is full and  Write wr_en flag is full is not asserted  
					 if (full_reg) NextState <= S4;
            	 else NextState <= S1;
            end	
				default: begin 
					 NextState <= S0;
            end				
		endcase
	end
	
	
	// L�gica combinacional de salida ************************************	
	always @* begin
	    case(State)
	        S0: begin  // Wait for start providing for initialization module
                reset_output_register <= 1'b1;
					 wr_en_reg <= 1'b0;
					 reset_file_register <= 1'b1;
					 enable_output_register <= 1'b0;
				end
				S1: begin // Wait for tlast
                reset_output_register <= 1'b1;
					 wr_en_reg <= 1'b0;
					 reset_file_register <= 1'b0;
					 enable_output_register <= 1'b0;
				end
				S2: begin // Wait for the last write in the file register
					 reset_output_register <= 1'b0;
					 wr_en_reg <= 1'b0;
					 reset_file_register <= 1'b0;
					 enable_output_register <= 1'b0;
				end
				S3: begin // Load output register and reset all the register file and counter
					 reset_output_register <= 1'b0;
					 wr_en_reg <= 1'b0;
					 reset_file_register <= 1'b1;
					 enable_output_register <= 1'b1;
            end	
				S4: begin // Wait if fifo is full and  Write wr_en flag is full is not asserted  
					 reset_output_register <= 1'b0;
					 if (full_reg) wr_en_reg <= 1'b0;
            	 else wr_en_reg <= 1'b1;
					 reset_file_register <= 1'b0;
					 enable_output_register <= 1'b0;
            end	
				default: begin 
					 reset_output_register <= 1'b1;
					 wr_en_reg <= 1'b0;
					 reset_file_register <= 1'b1;
					 enable_output_register <= 1'b0;
            end				
		endcase
	end
	
	// ******************************************************  ROM Memory ******************************************
	
	ROM ROM_BS_UID(user_clk, din_reg[(PACKET_SIZE-1-32):(PACKET_SIZE-1-32-7)] , BS_ID);
	
	// ******************************************************  Output register **************************************
	
	register #(.WIDTH(PACKET_SIZE)) Parallel_Output_Register (
		.user_clk(user_clk), 
		.RST(RST | reset_output_register), 
		.Enable(enable_output_register), 
		.D( {BS_ID, din_reg[PACKET_SIZE-1-8:0]} ), 
		.Q(din)
	);
	
	
	// **************************************** Error handler
	
	
   
   always @(posedge user_clk)
      if (RST)
         Q_seq_counter <= 0;
      else if (enable_output_register)
         Q_seq_counter <= Q_seq_counter + 1'b1;
	

   always @(posedge user_clk)
		if (RST) begin
			Error <= 1'b0;
		end else if (Enable_Registers[1]) begin
			if (Q_seq_counter == din_reg[PACKET_SIZE-1:PACKET_SIZE-8])
				Error <= 1'b0;
			else
				Error <= 1'b1;
	   end
	
	
	

endmodule



